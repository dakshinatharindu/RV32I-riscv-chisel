module ControlUnit(
  input  [31:0] io_instr,
  input         io_eq,
  input         io_ge,
  input         io_geu,
  input         io_valid,
  output [2:0]  io_format,
  output [3:0]  io_ALUCtrl,
  output        io_regWrite,
  output        io_memWrite,
  output        io_memRead,
  output        io_rs2Imm,
  output        io_aluMem,
  output        io_pcAluMem,
  output        io_pcImm,
  output        io_immBranch,
  output        io_aluBranch,
  output        io_stall,
  output [1:0]  io_storeType
);
  wire [6:0] opcode = io_instr[6:0]; // @[ControlUnit.scala 30:24]
  wire [6:0] func7 = io_instr[31:25]; // @[ControlUnit.scala 31:23]
  wire [2:0] func3 = io_instr[14:12]; // @[ControlUnit.scala 32:23]
  wire [4:0] subFormat = opcode[6:2]; // @[ControlUnit.scala 33:25]
  wire [3:0] funcCode = {func7[5],func3}; // @[ControlUnit.scala 34:27]
  wire [3:0] _GEN_1 = 4'h6 == funcCode ? 4'h1 : 4'h0; // @[ControlUnit.scala 62:24 71:28]
  wire [3:0] _GEN_2 = 4'hd == funcCode ? 4'h9 : _GEN_1; // @[ControlUnit.scala 62:24 70:29]
  wire [3:0] _GEN_3 = 4'h5 == funcCode ? 4'h8 : _GEN_2; // @[ControlUnit.scala 62:24 69:29]
  wire [3:0] _GEN_4 = 4'h4 == funcCode ? 4'h2 : _GEN_3; // @[ControlUnit.scala 62:24 68:29]
  wire [3:0] _GEN_5 = 4'h3 == funcCode ? 4'h7 : _GEN_4; // @[ControlUnit.scala 62:24 67:30]
  wire [3:0] _GEN_6 = 4'h2 == funcCode ? 4'h5 : _GEN_5; // @[ControlUnit.scala 62:24 66:29]
  wire [3:0] _GEN_7 = 4'h1 == funcCode ? 4'h6 : _GEN_6; // @[ControlUnit.scala 62:24 65:29]
  wire [3:0] _GEN_8 = 4'h8 == funcCode ? 4'h4 : _GEN_7; // @[ControlUnit.scala 62:24 64:29]
  wire [3:0] _GEN_9 = 4'h0 == funcCode ? 4'h3 : _GEN_8; // @[ControlUnit.scala 62:24 63:29]
  wire [3:0] _GEN_10 = ~funcCode[3] ? 4'h8 : 4'h9; // @[ControlUnit.scala 100:21 102:21 99:37]
  wire [3:0] _GEN_11 = 3'h5 == funcCode[2:0] ? _GEN_10 : 4'h0; // @[ControlUnit.scala 36:28 90:30]
  wire [3:0] _GEN_12 = 3'h1 == funcCode[2:0] ? 4'h6 : _GEN_11; // @[ControlUnit.scala 90:30 97:32]
  wire [3:0] _GEN_13 = 3'h7 == funcCode[2:0] ? 4'h0 : _GEN_12; // @[ControlUnit.scala 90:30 96:32]
  wire [3:0] _GEN_14 = 3'h6 == funcCode[2:0] ? 4'h1 : _GEN_13; // @[ControlUnit.scala 90:30 95:32]
  wire [3:0] _GEN_15 = 3'h4 == funcCode[2:0] ? 4'h2 : _GEN_14; // @[ControlUnit.scala 90:30 94:32]
  wire [3:0] _GEN_16 = 3'h3 == funcCode[2:0] ? 4'h7 : _GEN_15; // @[ControlUnit.scala 90:30 93:32]
  wire [3:0] _GEN_17 = 3'h2 == funcCode[2:0] ? 4'h5 : _GEN_16; // @[ControlUnit.scala 90:30 92:32]
  wire [3:0] _GEN_18 = 3'h0 == funcCode[2:0] ? 4'h3 : _GEN_17; // @[ControlUnit.scala 90:30 91:32]
  wire  _immBranch_T_1 = io_eq ? 1'h0 : 1'h1; // @[ControlUnit.scala 161:37]
  wire  _immBranch_T_2 = io_ge ? 1'h0 : 1'h1; // @[ControlUnit.scala 162:37]
  wire  _immBranch_T_4 = io_geu ? 1'h0 : 1'h1; // @[ControlUnit.scala 164:38]
  wire  _GEN_19 = 3'h7 == func3 & io_geu; // @[ControlUnit.scala 159:21 165:32 45:30]
  wire  _GEN_20 = 3'h6 == func3 ? _immBranch_T_4 : _GEN_19; // @[ControlUnit.scala 159:21 164:32]
  wire  _GEN_21 = 3'h5 == func3 ? io_ge : _GEN_20; // @[ControlUnit.scala 159:21 163:31]
  wire  _GEN_22 = 3'h4 == func3 ? _immBranch_T_2 : _GEN_21; // @[ControlUnit.scala 159:21 162:31]
  wire  _GEN_23 = 3'h1 == func3 ? _immBranch_T_1 : _GEN_22; // @[ControlUnit.scala 159:21 161:31]
  wire  _GEN_24 = 3'h0 == func3 ? io_eq : _GEN_23; // @[ControlUnit.scala 159:21 160:31]
  wire [2:0] _GEN_27 = 5'h1b == subFormat ? 3'h5 : 3'h0; // @[ControlUnit.scala 218:14 49:21 37:27]
  wire  _GEN_30 = 5'h5 == subFormat ? 1'h0 : 5'h1b == subFormat; // @[ControlUnit.scala 197:17 49:21]
  wire  _GEN_31 = 5'h5 == subFormat | 5'h1b == subFormat; // @[ControlUnit.scala 199:13 49:21]
  wire [2:0] _GEN_32 = 5'h5 == subFormat ? 3'h4 : _GEN_27; // @[ControlUnit.scala 205:14 49:21]
  wire  _GEN_35 = 5'hd == subFormat ? 1'h0 : _GEN_30; // @[ControlUnit.scala 181:17 49:21]
  wire  _GEN_37 = 5'hd == subFormat | _GEN_31; // @[ControlUnit.scala 183:13 49:21]
  wire [3:0] _GEN_38 = 5'hd == subFormat ? 4'hb : 4'h0; // @[ControlUnit.scala 189:15 49:21 36:28]
  wire [2:0] _GEN_39 = 5'hd == subFormat ? 3'h4 : _GEN_32; // @[ControlUnit.scala 191:14 49:21]
  wire  _GEN_40 = 5'hd == subFormat ? 1'h0 : 5'h5 == subFormat; // @[ControlUnit.scala 49:21 44:26]
  wire  _GEN_42 = 5'h18 == subFormat ? _GEN_24 : _GEN_35; // @[ControlUnit.scala 49:21]
  wire  _GEN_44 = 5'h18 == subFormat | _GEN_37; // @[ControlUnit.scala 168:13 49:21]
  wire  _GEN_45 = 5'h18 == subFormat ? 1'h0 : _GEN_37; // @[ControlUnit.scala 170:16 49:21]
  wire [2:0] _GEN_46 = 5'h18 == subFormat ? 3'h3 : _GEN_39; // @[ControlUnit.scala 174:14 49:21]
  wire  _GEN_47 = 5'h18 == subFormat ? 1'h0 : 5'hd == subFormat; // @[ControlUnit.scala 49:21 43:29]
  wire [3:0] _GEN_48 = 5'h18 == subFormat ? 4'h0 : _GEN_38; // @[ControlUnit.scala 49:21 36:28]
  wire  _GEN_49 = 5'h18 == subFormat ? 1'h0 : _GEN_40; // @[ControlUnit.scala 49:21 44:26]
  wire  _GEN_51 = 5'h8 == subFormat ? 1'h0 : _GEN_42; // @[ControlUnit.scala 144:17 49:21]
  wire  _GEN_53 = 5'h8 == subFormat ? io_valid : _GEN_44; // @[ControlUnit.scala 146:13 49:21]
  wire  _GEN_54 = 5'h8 == subFormat ? 1'h0 : _GEN_45; // @[ControlUnit.scala 148:16 49:21]
  wire [3:0] _GEN_56 = 5'h8 == subFormat ? 4'h3 : _GEN_48; // @[ControlUnit.scala 152:15 49:21]
  wire [2:0] _GEN_57 = 5'h8 == subFormat ? 3'h2 : _GEN_46; // @[ControlUnit.scala 154:14 49:21]
  wire  _GEN_59 = 5'h8 == subFormat ? 1'h0 : _GEN_47; // @[ControlUnit.scala 49:21 43:29]
  wire  _GEN_60 = 5'h8 == subFormat ? 1'h0 : _GEN_49; // @[ControlUnit.scala 49:21 44:26]
  wire  _GEN_61 = 5'h19 == subFormat ? 1'h0 : _GEN_60; // @[ControlUnit.scala 128:13 49:21]
  wire  _GEN_62 = 5'h19 == subFormat ? 1'h0 : _GEN_59; // @[ControlUnit.scala 129:16 49:21]
  wire  _GEN_64 = 5'h19 == subFormat | _GEN_53; // @[ControlUnit.scala 131:13 49:21]
  wire  _GEN_65 = 5'h19 == subFormat | _GEN_54; // @[ControlUnit.scala 133:16 49:21]
  wire  _GEN_67 = 5'h19 == subFormat ? 1'h0 : 5'h8 == subFormat; // @[ControlUnit.scala 135:16 49:21]
  wire [3:0] _GEN_68 = 5'h19 == subFormat ? 4'ha : _GEN_56; // @[ControlUnit.scala 137:15 49:21]
  wire [2:0] _GEN_69 = 5'h19 == subFormat ? 3'h1 : _GEN_57; // @[ControlUnit.scala 139:14 49:21]
  wire  _GEN_71 = 5'h19 == subFormat ? 1'h0 : _GEN_51; // @[ControlUnit.scala 49:21 45:30]
  wire  _GEN_73 = 5'h0 == subFormat | _GEN_67; // @[ControlUnit.scala 111:14 49:21]
  wire  _GEN_75 = 5'h0 == subFormat | _GEN_62; // @[ControlUnit.scala 113:16 49:21]
  wire  _GEN_76 = 5'h0 == subFormat ? 1'h0 : _GEN_71; // @[ControlUnit.scala 114:17 49:21]
  wire  _GEN_77 = 5'h0 == subFormat ? 1'h0 : 5'h19 == subFormat; // @[ControlUnit.scala 115:17 49:21]
  wire  _GEN_78 = 5'h0 == subFormat ? io_valid : _GEN_64; // @[ControlUnit.scala 116:13 49:21]
  wire  _GEN_79 = 5'h0 == subFormat | _GEN_65; // @[ControlUnit.scala 118:16 49:21]
  wire  _GEN_81 = 5'h0 == subFormat ? 1'h0 : _GEN_67; // @[ControlUnit.scala 120:16 49:21]
  wire [3:0] _GEN_82 = 5'h0 == subFormat ? 4'h3 : _GEN_68; // @[ControlUnit.scala 122:15 49:21]
  wire [2:0] _GEN_83 = 5'h0 == subFormat ? 3'h1 : _GEN_69; // @[ControlUnit.scala 124:14 49:21]
  wire  _GEN_84 = 5'h0 == subFormat ? 1'h0 : _GEN_61; // @[ControlUnit.scala 49:21 44:26]
  wire  _GEN_85 = 5'h4 == subFormat | _GEN_73; // @[ControlUnit.scala 49:21 79:14]
  wire  _GEN_86 = 5'h4 == subFormat ? 1'h0 : 5'h0 == subFormat; // @[ControlUnit.scala 49:21 80:14]
  wire  _GEN_87 = 5'h4 == subFormat | _GEN_75; // @[ControlUnit.scala 49:21 81:16]
  wire  _GEN_88 = 5'h4 == subFormat ? 1'h0 : _GEN_76; // @[ControlUnit.scala 49:21 82:17]
  wire  _GEN_89 = 5'h4 == subFormat ? 1'h0 : _GEN_77; // @[ControlUnit.scala 49:21 83:17]
  wire  _GEN_90 = 5'h4 == subFormat | _GEN_78; // @[ControlUnit.scala 49:21 84:13]
  wire  _GEN_91 = 5'h4 == subFormat | _GEN_79; // @[ControlUnit.scala 49:21 86:16]
  wire  _GEN_93 = 5'h4 == subFormat ? 1'h0 : _GEN_81; // @[ControlUnit.scala 49:21 88:16]
  wire [3:0] _GEN_94 = 5'h4 == subFormat ? _GEN_18 : _GEN_82; // @[ControlUnit.scala 49:21]
  wire [2:0] _GEN_95 = 5'h4 == subFormat ? 3'h1 : _GEN_83; // @[ControlUnit.scala 107:14 49:21]
  wire  _GEN_96 = 5'h4 == subFormat ? 1'h0 : _GEN_84; // @[ControlUnit.scala 49:21 44:26]
  assign io_format = 5'hc == subFormat ? 3'h0 : _GEN_95; // @[ControlUnit.scala 49:21 75:14]
  assign io_ALUCtrl = 5'hc == subFormat ? _GEN_9 : _GEN_94; // @[ControlUnit.scala 49:21]
  assign io_regWrite = 5'hc == subFormat | _GEN_91; // @[ControlUnit.scala 49:21 58:16]
  assign io_memWrite = 5'hc == subFormat ? 1'h0 : _GEN_93; // @[ControlUnit.scala 49:21 60:16]
  assign io_memRead = 5'hc == subFormat ? 1'h0 : _GEN_86; // @[ControlUnit.scala 49:21 59:15]
  assign io_rs2Imm = 5'hc == subFormat ? 1'h0 : _GEN_85; // @[ControlUnit.scala 49:21 51:14]
  assign io_aluMem = 5'hc == subFormat ? 1'h0 : _GEN_86; // @[ControlUnit.scala 49:21 52:14]
  assign io_pcAluMem = 5'hc == subFormat | _GEN_87; // @[ControlUnit.scala 49:21 53:16]
  assign io_pcImm = 5'hc == subFormat ? 1'h0 : _GEN_96; // @[ControlUnit.scala 49:21 44:26]
  assign io_immBranch = 5'hc == subFormat ? 1'h0 : _GEN_88; // @[ControlUnit.scala 49:21 54:17]
  assign io_aluBranch = 5'hc == subFormat ? 1'h0 : _GEN_89; // @[ControlUnit.scala 49:21 55:17]
  assign io_stall = 5'hc == subFormat | _GEN_90; // @[ControlUnit.scala 49:21 56:13]
  assign io_storeType = func3[1:0]; // @[ControlUnit.scala 234:24]
endmodule
module RegisterFile(
  input         clock,
  input         reset,
  input  [4:0]  io_readAddr1,
  input  [4:0]  io_readAddr2,
  input  [4:0]  io_writeAddr,
  input  [31:0] io_writeData,
  input         io_writeEn,
  output [31:0] io_readData1,
  output [31:0] io_readData2
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] registerFile_0; // @[RegisterFile.scala 19:29]
  reg [31:0] registerFile_1; // @[RegisterFile.scala 19:29]
  reg [31:0] registerFile_2; // @[RegisterFile.scala 19:29]
  reg [31:0] registerFile_3; // @[RegisterFile.scala 19:29]
  reg [31:0] registerFile_4; // @[RegisterFile.scala 19:29]
  reg [31:0] registerFile_5; // @[RegisterFile.scala 19:29]
  reg [31:0] registerFile_6; // @[RegisterFile.scala 19:29]
  reg [31:0] registerFile_7; // @[RegisterFile.scala 19:29]
  reg [31:0] registerFile_8; // @[RegisterFile.scala 19:29]
  reg [31:0] registerFile_9; // @[RegisterFile.scala 19:29]
  reg [31:0] registerFile_10; // @[RegisterFile.scala 19:29]
  reg [31:0] registerFile_11; // @[RegisterFile.scala 19:29]
  reg [31:0] registerFile_12; // @[RegisterFile.scala 19:29]
  reg [31:0] registerFile_13; // @[RegisterFile.scala 19:29]
  reg [31:0] registerFile_14; // @[RegisterFile.scala 19:29]
  reg [31:0] registerFile_15; // @[RegisterFile.scala 19:29]
  reg [31:0] registerFile_16; // @[RegisterFile.scala 19:29]
  reg [31:0] registerFile_17; // @[RegisterFile.scala 19:29]
  reg [31:0] registerFile_18; // @[RegisterFile.scala 19:29]
  reg [31:0] registerFile_19; // @[RegisterFile.scala 19:29]
  reg [31:0] registerFile_20; // @[RegisterFile.scala 19:29]
  reg [31:0] registerFile_21; // @[RegisterFile.scala 19:29]
  reg [31:0] registerFile_22; // @[RegisterFile.scala 19:29]
  reg [31:0] registerFile_23; // @[RegisterFile.scala 19:29]
  reg [31:0] registerFile_24; // @[RegisterFile.scala 19:29]
  reg [31:0] registerFile_25; // @[RegisterFile.scala 19:29]
  reg [31:0] registerFile_26; // @[RegisterFile.scala 19:29]
  reg [31:0] registerFile_27; // @[RegisterFile.scala 19:29]
  reg [31:0] registerFile_28; // @[RegisterFile.scala 19:29]
  reg [31:0] registerFile_29; // @[RegisterFile.scala 19:29]
  reg [31:0] registerFile_30; // @[RegisterFile.scala 19:29]
  reg [31:0] registerFile_31; // @[RegisterFile.scala 19:29]
  wire [31:0] _GEN_1 = 5'h1 == io_readAddr1 ? $signed(registerFile_1) : $signed(registerFile_0); // @[RegisterFile.scala 23:{18,18}]
  wire [31:0] _GEN_2 = 5'h2 == io_readAddr1 ? $signed(registerFile_2) : $signed(_GEN_1); // @[RegisterFile.scala 23:{18,18}]
  wire [31:0] _GEN_3 = 5'h3 == io_readAddr1 ? $signed(registerFile_3) : $signed(_GEN_2); // @[RegisterFile.scala 23:{18,18}]
  wire [31:0] _GEN_4 = 5'h4 == io_readAddr1 ? $signed(registerFile_4) : $signed(_GEN_3); // @[RegisterFile.scala 23:{18,18}]
  wire [31:0] _GEN_5 = 5'h5 == io_readAddr1 ? $signed(registerFile_5) : $signed(_GEN_4); // @[RegisterFile.scala 23:{18,18}]
  wire [31:0] _GEN_6 = 5'h6 == io_readAddr1 ? $signed(registerFile_6) : $signed(_GEN_5); // @[RegisterFile.scala 23:{18,18}]
  wire [31:0] _GEN_7 = 5'h7 == io_readAddr1 ? $signed(registerFile_7) : $signed(_GEN_6); // @[RegisterFile.scala 23:{18,18}]
  wire [31:0] _GEN_8 = 5'h8 == io_readAddr1 ? $signed(registerFile_8) : $signed(_GEN_7); // @[RegisterFile.scala 23:{18,18}]
  wire [31:0] _GEN_9 = 5'h9 == io_readAddr1 ? $signed(registerFile_9) : $signed(_GEN_8); // @[RegisterFile.scala 23:{18,18}]
  wire [31:0] _GEN_10 = 5'ha == io_readAddr1 ? $signed(registerFile_10) : $signed(_GEN_9); // @[RegisterFile.scala 23:{18,18}]
  wire [31:0] _GEN_11 = 5'hb == io_readAddr1 ? $signed(registerFile_11) : $signed(_GEN_10); // @[RegisterFile.scala 23:{18,18}]
  wire [31:0] _GEN_12 = 5'hc == io_readAddr1 ? $signed(registerFile_12) : $signed(_GEN_11); // @[RegisterFile.scala 23:{18,18}]
  wire [31:0] _GEN_13 = 5'hd == io_readAddr1 ? $signed(registerFile_13) : $signed(_GEN_12); // @[RegisterFile.scala 23:{18,18}]
  wire [31:0] _GEN_14 = 5'he == io_readAddr1 ? $signed(registerFile_14) : $signed(_GEN_13); // @[RegisterFile.scala 23:{18,18}]
  wire [31:0] _GEN_15 = 5'hf == io_readAddr1 ? $signed(registerFile_15) : $signed(_GEN_14); // @[RegisterFile.scala 23:{18,18}]
  wire [31:0] _GEN_16 = 5'h10 == io_readAddr1 ? $signed(registerFile_16) : $signed(_GEN_15); // @[RegisterFile.scala 23:{18,18}]
  wire [31:0] _GEN_17 = 5'h11 == io_readAddr1 ? $signed(registerFile_17) : $signed(_GEN_16); // @[RegisterFile.scala 23:{18,18}]
  wire [31:0] _GEN_18 = 5'h12 == io_readAddr1 ? $signed(registerFile_18) : $signed(_GEN_17); // @[RegisterFile.scala 23:{18,18}]
  wire [31:0] _GEN_19 = 5'h13 == io_readAddr1 ? $signed(registerFile_19) : $signed(_GEN_18); // @[RegisterFile.scala 23:{18,18}]
  wire [31:0] _GEN_20 = 5'h14 == io_readAddr1 ? $signed(registerFile_20) : $signed(_GEN_19); // @[RegisterFile.scala 23:{18,18}]
  wire [31:0] _GEN_21 = 5'h15 == io_readAddr1 ? $signed(registerFile_21) : $signed(_GEN_20); // @[RegisterFile.scala 23:{18,18}]
  wire [31:0] _GEN_22 = 5'h16 == io_readAddr1 ? $signed(registerFile_22) : $signed(_GEN_21); // @[RegisterFile.scala 23:{18,18}]
  wire [31:0] _GEN_23 = 5'h17 == io_readAddr1 ? $signed(registerFile_23) : $signed(_GEN_22); // @[RegisterFile.scala 23:{18,18}]
  wire [31:0] _GEN_24 = 5'h18 == io_readAddr1 ? $signed(registerFile_24) : $signed(_GEN_23); // @[RegisterFile.scala 23:{18,18}]
  wire [31:0] _GEN_25 = 5'h19 == io_readAddr1 ? $signed(registerFile_25) : $signed(_GEN_24); // @[RegisterFile.scala 23:{18,18}]
  wire [31:0] _GEN_26 = 5'h1a == io_readAddr1 ? $signed(registerFile_26) : $signed(_GEN_25); // @[RegisterFile.scala 23:{18,18}]
  wire [31:0] _GEN_27 = 5'h1b == io_readAddr1 ? $signed(registerFile_27) : $signed(_GEN_26); // @[RegisterFile.scala 23:{18,18}]
  wire [31:0] _GEN_28 = 5'h1c == io_readAddr1 ? $signed(registerFile_28) : $signed(_GEN_27); // @[RegisterFile.scala 23:{18,18}]
  wire [31:0] _GEN_29 = 5'h1d == io_readAddr1 ? $signed(registerFile_29) : $signed(_GEN_28); // @[RegisterFile.scala 23:{18,18}]
  wire [31:0] _GEN_30 = 5'h1e == io_readAddr1 ? $signed(registerFile_30) : $signed(_GEN_29); // @[RegisterFile.scala 23:{18,18}]
  wire [31:0] _GEN_31 = 5'h1f == io_readAddr1 ? $signed(registerFile_31) : $signed(_GEN_30); // @[RegisterFile.scala 23:{18,18}]
  wire [31:0] _GEN_34 = 5'h1 == io_readAddr2 ? $signed(registerFile_1) : $signed(registerFile_0); // @[RegisterFile.scala 29:{18,18}]
  wire [31:0] _GEN_35 = 5'h2 == io_readAddr2 ? $signed(registerFile_2) : $signed(_GEN_34); // @[RegisterFile.scala 29:{18,18}]
  wire [31:0] _GEN_36 = 5'h3 == io_readAddr2 ? $signed(registerFile_3) : $signed(_GEN_35); // @[RegisterFile.scala 29:{18,18}]
  wire [31:0] _GEN_37 = 5'h4 == io_readAddr2 ? $signed(registerFile_4) : $signed(_GEN_36); // @[RegisterFile.scala 29:{18,18}]
  wire [31:0] _GEN_38 = 5'h5 == io_readAddr2 ? $signed(registerFile_5) : $signed(_GEN_37); // @[RegisterFile.scala 29:{18,18}]
  wire [31:0] _GEN_39 = 5'h6 == io_readAddr2 ? $signed(registerFile_6) : $signed(_GEN_38); // @[RegisterFile.scala 29:{18,18}]
  wire [31:0] _GEN_40 = 5'h7 == io_readAddr2 ? $signed(registerFile_7) : $signed(_GEN_39); // @[RegisterFile.scala 29:{18,18}]
  wire [31:0] _GEN_41 = 5'h8 == io_readAddr2 ? $signed(registerFile_8) : $signed(_GEN_40); // @[RegisterFile.scala 29:{18,18}]
  wire [31:0] _GEN_42 = 5'h9 == io_readAddr2 ? $signed(registerFile_9) : $signed(_GEN_41); // @[RegisterFile.scala 29:{18,18}]
  wire [31:0] _GEN_43 = 5'ha == io_readAddr2 ? $signed(registerFile_10) : $signed(_GEN_42); // @[RegisterFile.scala 29:{18,18}]
  wire [31:0] _GEN_44 = 5'hb == io_readAddr2 ? $signed(registerFile_11) : $signed(_GEN_43); // @[RegisterFile.scala 29:{18,18}]
  wire [31:0] _GEN_45 = 5'hc == io_readAddr2 ? $signed(registerFile_12) : $signed(_GEN_44); // @[RegisterFile.scala 29:{18,18}]
  wire [31:0] _GEN_46 = 5'hd == io_readAddr2 ? $signed(registerFile_13) : $signed(_GEN_45); // @[RegisterFile.scala 29:{18,18}]
  wire [31:0] _GEN_47 = 5'he == io_readAddr2 ? $signed(registerFile_14) : $signed(_GEN_46); // @[RegisterFile.scala 29:{18,18}]
  wire [31:0] _GEN_48 = 5'hf == io_readAddr2 ? $signed(registerFile_15) : $signed(_GEN_47); // @[RegisterFile.scala 29:{18,18}]
  wire [31:0] _GEN_49 = 5'h10 == io_readAddr2 ? $signed(registerFile_16) : $signed(_GEN_48); // @[RegisterFile.scala 29:{18,18}]
  wire [31:0] _GEN_50 = 5'h11 == io_readAddr2 ? $signed(registerFile_17) : $signed(_GEN_49); // @[RegisterFile.scala 29:{18,18}]
  wire [31:0] _GEN_51 = 5'h12 == io_readAddr2 ? $signed(registerFile_18) : $signed(_GEN_50); // @[RegisterFile.scala 29:{18,18}]
  wire [31:0] _GEN_52 = 5'h13 == io_readAddr2 ? $signed(registerFile_19) : $signed(_GEN_51); // @[RegisterFile.scala 29:{18,18}]
  wire [31:0] _GEN_53 = 5'h14 == io_readAddr2 ? $signed(registerFile_20) : $signed(_GEN_52); // @[RegisterFile.scala 29:{18,18}]
  wire [31:0] _GEN_54 = 5'h15 == io_readAddr2 ? $signed(registerFile_21) : $signed(_GEN_53); // @[RegisterFile.scala 29:{18,18}]
  wire [31:0] _GEN_55 = 5'h16 == io_readAddr2 ? $signed(registerFile_22) : $signed(_GEN_54); // @[RegisterFile.scala 29:{18,18}]
  wire [31:0] _GEN_56 = 5'h17 == io_readAddr2 ? $signed(registerFile_23) : $signed(_GEN_55); // @[RegisterFile.scala 29:{18,18}]
  wire [31:0] _GEN_57 = 5'h18 == io_readAddr2 ? $signed(registerFile_24) : $signed(_GEN_56); // @[RegisterFile.scala 29:{18,18}]
  wire [31:0] _GEN_58 = 5'h19 == io_readAddr2 ? $signed(registerFile_25) : $signed(_GEN_57); // @[RegisterFile.scala 29:{18,18}]
  wire [31:0] _GEN_59 = 5'h1a == io_readAddr2 ? $signed(registerFile_26) : $signed(_GEN_58); // @[RegisterFile.scala 29:{18,18}]
  wire [31:0] _GEN_60 = 5'h1b == io_readAddr2 ? $signed(registerFile_27) : $signed(_GEN_59); // @[RegisterFile.scala 29:{18,18}]
  wire [31:0] _GEN_61 = 5'h1c == io_readAddr2 ? $signed(registerFile_28) : $signed(_GEN_60); // @[RegisterFile.scala 29:{18,18}]
  wire [31:0] _GEN_62 = 5'h1d == io_readAddr2 ? $signed(registerFile_29) : $signed(_GEN_61); // @[RegisterFile.scala 29:{18,18}]
  wire [31:0] _GEN_63 = 5'h1e == io_readAddr2 ? $signed(registerFile_30) : $signed(_GEN_62); // @[RegisterFile.scala 29:{18,18}]
  wire [31:0] _GEN_64 = 5'h1f == io_readAddr2 ? $signed(registerFile_31) : $signed(_GEN_63); // @[RegisterFile.scala 29:{18,18}]
  assign io_readData1 = io_readAddr1 == 5'h0 ? $signed(32'sh0) : $signed(_GEN_31); // @[RegisterFile.scala 20:30 21:18 23:18]
  assign io_readData2 = io_readAddr2 == 5'h0 ? $signed(32'sh0) : $signed(_GEN_64); // @[RegisterFile.scala 26:30 27:18 29:18]
  always @(posedge clock) begin
    if (reset) begin // @[RegisterFile.scala 19:29]
      registerFile_0 <= 32'sh0; // @[RegisterFile.scala 19:29]
    end else if (io_writeEn) begin // @[RegisterFile.scala 32:20]
      if (5'h0 == io_writeAddr) begin // @[RegisterFile.scala 33:32]
        registerFile_0 <= io_writeData; // @[RegisterFile.scala 33:32]
      end
    end
    if (reset) begin // @[RegisterFile.scala 19:29]
      registerFile_1 <= 32'sh0; // @[RegisterFile.scala 19:29]
    end else if (io_writeEn) begin // @[RegisterFile.scala 32:20]
      if (5'h1 == io_writeAddr) begin // @[RegisterFile.scala 33:32]
        registerFile_1 <= io_writeData; // @[RegisterFile.scala 33:32]
      end
    end
    if (reset) begin // @[RegisterFile.scala 19:29]
      registerFile_2 <= 32'sh0; // @[RegisterFile.scala 19:29]
    end else if (io_writeEn) begin // @[RegisterFile.scala 32:20]
      if (5'h2 == io_writeAddr) begin // @[RegisterFile.scala 33:32]
        registerFile_2 <= io_writeData; // @[RegisterFile.scala 33:32]
      end
    end
    if (reset) begin // @[RegisterFile.scala 19:29]
      registerFile_3 <= 32'sh0; // @[RegisterFile.scala 19:29]
    end else if (io_writeEn) begin // @[RegisterFile.scala 32:20]
      if (5'h3 == io_writeAddr) begin // @[RegisterFile.scala 33:32]
        registerFile_3 <= io_writeData; // @[RegisterFile.scala 33:32]
      end
    end
    if (reset) begin // @[RegisterFile.scala 19:29]
      registerFile_4 <= 32'sh0; // @[RegisterFile.scala 19:29]
    end else if (io_writeEn) begin // @[RegisterFile.scala 32:20]
      if (5'h4 == io_writeAddr) begin // @[RegisterFile.scala 33:32]
        registerFile_4 <= io_writeData; // @[RegisterFile.scala 33:32]
      end
    end
    if (reset) begin // @[RegisterFile.scala 19:29]
      registerFile_5 <= 32'sh0; // @[RegisterFile.scala 19:29]
    end else if (io_writeEn) begin // @[RegisterFile.scala 32:20]
      if (5'h5 == io_writeAddr) begin // @[RegisterFile.scala 33:32]
        registerFile_5 <= io_writeData; // @[RegisterFile.scala 33:32]
      end
    end
    if (reset) begin // @[RegisterFile.scala 19:29]
      registerFile_6 <= 32'sh0; // @[RegisterFile.scala 19:29]
    end else if (io_writeEn) begin // @[RegisterFile.scala 32:20]
      if (5'h6 == io_writeAddr) begin // @[RegisterFile.scala 33:32]
        registerFile_6 <= io_writeData; // @[RegisterFile.scala 33:32]
      end
    end
    if (reset) begin // @[RegisterFile.scala 19:29]
      registerFile_7 <= 32'sh0; // @[RegisterFile.scala 19:29]
    end else if (io_writeEn) begin // @[RegisterFile.scala 32:20]
      if (5'h7 == io_writeAddr) begin // @[RegisterFile.scala 33:32]
        registerFile_7 <= io_writeData; // @[RegisterFile.scala 33:32]
      end
    end
    if (reset) begin // @[RegisterFile.scala 19:29]
      registerFile_8 <= 32'sh0; // @[RegisterFile.scala 19:29]
    end else if (io_writeEn) begin // @[RegisterFile.scala 32:20]
      if (5'h8 == io_writeAddr) begin // @[RegisterFile.scala 33:32]
        registerFile_8 <= io_writeData; // @[RegisterFile.scala 33:32]
      end
    end
    if (reset) begin // @[RegisterFile.scala 19:29]
      registerFile_9 <= 32'sh0; // @[RegisterFile.scala 19:29]
    end else if (io_writeEn) begin // @[RegisterFile.scala 32:20]
      if (5'h9 == io_writeAddr) begin // @[RegisterFile.scala 33:32]
        registerFile_9 <= io_writeData; // @[RegisterFile.scala 33:32]
      end
    end
    if (reset) begin // @[RegisterFile.scala 19:29]
      registerFile_10 <= 32'sh0; // @[RegisterFile.scala 19:29]
    end else if (io_writeEn) begin // @[RegisterFile.scala 32:20]
      if (5'ha == io_writeAddr) begin // @[RegisterFile.scala 33:32]
        registerFile_10 <= io_writeData; // @[RegisterFile.scala 33:32]
      end
    end
    if (reset) begin // @[RegisterFile.scala 19:29]
      registerFile_11 <= 32'sh0; // @[RegisterFile.scala 19:29]
    end else if (io_writeEn) begin // @[RegisterFile.scala 32:20]
      if (5'hb == io_writeAddr) begin // @[RegisterFile.scala 33:32]
        registerFile_11 <= io_writeData; // @[RegisterFile.scala 33:32]
      end
    end
    if (reset) begin // @[RegisterFile.scala 19:29]
      registerFile_12 <= 32'sh0; // @[RegisterFile.scala 19:29]
    end else if (io_writeEn) begin // @[RegisterFile.scala 32:20]
      if (5'hc == io_writeAddr) begin // @[RegisterFile.scala 33:32]
        registerFile_12 <= io_writeData; // @[RegisterFile.scala 33:32]
      end
    end
    if (reset) begin // @[RegisterFile.scala 19:29]
      registerFile_13 <= 32'sh0; // @[RegisterFile.scala 19:29]
    end else if (io_writeEn) begin // @[RegisterFile.scala 32:20]
      if (5'hd == io_writeAddr) begin // @[RegisterFile.scala 33:32]
        registerFile_13 <= io_writeData; // @[RegisterFile.scala 33:32]
      end
    end
    if (reset) begin // @[RegisterFile.scala 19:29]
      registerFile_14 <= 32'sh0; // @[RegisterFile.scala 19:29]
    end else if (io_writeEn) begin // @[RegisterFile.scala 32:20]
      if (5'he == io_writeAddr) begin // @[RegisterFile.scala 33:32]
        registerFile_14 <= io_writeData; // @[RegisterFile.scala 33:32]
      end
    end
    if (reset) begin // @[RegisterFile.scala 19:29]
      registerFile_15 <= 32'sh0; // @[RegisterFile.scala 19:29]
    end else if (io_writeEn) begin // @[RegisterFile.scala 32:20]
      if (5'hf == io_writeAddr) begin // @[RegisterFile.scala 33:32]
        registerFile_15 <= io_writeData; // @[RegisterFile.scala 33:32]
      end
    end
    if (reset) begin // @[RegisterFile.scala 19:29]
      registerFile_16 <= 32'sh0; // @[RegisterFile.scala 19:29]
    end else if (io_writeEn) begin // @[RegisterFile.scala 32:20]
      if (5'h10 == io_writeAddr) begin // @[RegisterFile.scala 33:32]
        registerFile_16 <= io_writeData; // @[RegisterFile.scala 33:32]
      end
    end
    if (reset) begin // @[RegisterFile.scala 19:29]
      registerFile_17 <= 32'sh0; // @[RegisterFile.scala 19:29]
    end else if (io_writeEn) begin // @[RegisterFile.scala 32:20]
      if (5'h11 == io_writeAddr) begin // @[RegisterFile.scala 33:32]
        registerFile_17 <= io_writeData; // @[RegisterFile.scala 33:32]
      end
    end
    if (reset) begin // @[RegisterFile.scala 19:29]
      registerFile_18 <= 32'sh0; // @[RegisterFile.scala 19:29]
    end else if (io_writeEn) begin // @[RegisterFile.scala 32:20]
      if (5'h12 == io_writeAddr) begin // @[RegisterFile.scala 33:32]
        registerFile_18 <= io_writeData; // @[RegisterFile.scala 33:32]
      end
    end
    if (reset) begin // @[RegisterFile.scala 19:29]
      registerFile_19 <= 32'sh0; // @[RegisterFile.scala 19:29]
    end else if (io_writeEn) begin // @[RegisterFile.scala 32:20]
      if (5'h13 == io_writeAddr) begin // @[RegisterFile.scala 33:32]
        registerFile_19 <= io_writeData; // @[RegisterFile.scala 33:32]
      end
    end
    if (reset) begin // @[RegisterFile.scala 19:29]
      registerFile_20 <= 32'sh0; // @[RegisterFile.scala 19:29]
    end else if (io_writeEn) begin // @[RegisterFile.scala 32:20]
      if (5'h14 == io_writeAddr) begin // @[RegisterFile.scala 33:32]
        registerFile_20 <= io_writeData; // @[RegisterFile.scala 33:32]
      end
    end
    if (reset) begin // @[RegisterFile.scala 19:29]
      registerFile_21 <= 32'sh0; // @[RegisterFile.scala 19:29]
    end else if (io_writeEn) begin // @[RegisterFile.scala 32:20]
      if (5'h15 == io_writeAddr) begin // @[RegisterFile.scala 33:32]
        registerFile_21 <= io_writeData; // @[RegisterFile.scala 33:32]
      end
    end
    if (reset) begin // @[RegisterFile.scala 19:29]
      registerFile_22 <= 32'sh0; // @[RegisterFile.scala 19:29]
    end else if (io_writeEn) begin // @[RegisterFile.scala 32:20]
      if (5'h16 == io_writeAddr) begin // @[RegisterFile.scala 33:32]
        registerFile_22 <= io_writeData; // @[RegisterFile.scala 33:32]
      end
    end
    if (reset) begin // @[RegisterFile.scala 19:29]
      registerFile_23 <= 32'sh0; // @[RegisterFile.scala 19:29]
    end else if (io_writeEn) begin // @[RegisterFile.scala 32:20]
      if (5'h17 == io_writeAddr) begin // @[RegisterFile.scala 33:32]
        registerFile_23 <= io_writeData; // @[RegisterFile.scala 33:32]
      end
    end
    if (reset) begin // @[RegisterFile.scala 19:29]
      registerFile_24 <= 32'sh0; // @[RegisterFile.scala 19:29]
    end else if (io_writeEn) begin // @[RegisterFile.scala 32:20]
      if (5'h18 == io_writeAddr) begin // @[RegisterFile.scala 33:32]
        registerFile_24 <= io_writeData; // @[RegisterFile.scala 33:32]
      end
    end
    if (reset) begin // @[RegisterFile.scala 19:29]
      registerFile_25 <= 32'sh0; // @[RegisterFile.scala 19:29]
    end else if (io_writeEn) begin // @[RegisterFile.scala 32:20]
      if (5'h19 == io_writeAddr) begin // @[RegisterFile.scala 33:32]
        registerFile_25 <= io_writeData; // @[RegisterFile.scala 33:32]
      end
    end
    if (reset) begin // @[RegisterFile.scala 19:29]
      registerFile_26 <= 32'sh0; // @[RegisterFile.scala 19:29]
    end else if (io_writeEn) begin // @[RegisterFile.scala 32:20]
      if (5'h1a == io_writeAddr) begin // @[RegisterFile.scala 33:32]
        registerFile_26 <= io_writeData; // @[RegisterFile.scala 33:32]
      end
    end
    if (reset) begin // @[RegisterFile.scala 19:29]
      registerFile_27 <= 32'sh0; // @[RegisterFile.scala 19:29]
    end else if (io_writeEn) begin // @[RegisterFile.scala 32:20]
      if (5'h1b == io_writeAddr) begin // @[RegisterFile.scala 33:32]
        registerFile_27 <= io_writeData; // @[RegisterFile.scala 33:32]
      end
    end
    if (reset) begin // @[RegisterFile.scala 19:29]
      registerFile_28 <= 32'sh0; // @[RegisterFile.scala 19:29]
    end else if (io_writeEn) begin // @[RegisterFile.scala 32:20]
      if (5'h1c == io_writeAddr) begin // @[RegisterFile.scala 33:32]
        registerFile_28 <= io_writeData; // @[RegisterFile.scala 33:32]
      end
    end
    if (reset) begin // @[RegisterFile.scala 19:29]
      registerFile_29 <= 32'sh0; // @[RegisterFile.scala 19:29]
    end else if (io_writeEn) begin // @[RegisterFile.scala 32:20]
      if (5'h1d == io_writeAddr) begin // @[RegisterFile.scala 33:32]
        registerFile_29 <= io_writeData; // @[RegisterFile.scala 33:32]
      end
    end
    if (reset) begin // @[RegisterFile.scala 19:29]
      registerFile_30 <= 32'sh0; // @[RegisterFile.scala 19:29]
    end else if (io_writeEn) begin // @[RegisterFile.scala 32:20]
      if (5'h1e == io_writeAddr) begin // @[RegisterFile.scala 33:32]
        registerFile_30 <= io_writeData; // @[RegisterFile.scala 33:32]
      end
    end
    if (reset) begin // @[RegisterFile.scala 19:29]
      registerFile_31 <= 32'sh0; // @[RegisterFile.scala 19:29]
    end else if (io_writeEn) begin // @[RegisterFile.scala 32:20]
      if (5'h1f == io_writeAddr) begin // @[RegisterFile.scala 33:32]
        registerFile_31 <= io_writeData; // @[RegisterFile.scala 33:32]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  registerFile_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  registerFile_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  registerFile_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  registerFile_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  registerFile_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  registerFile_5 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  registerFile_6 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  registerFile_7 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  registerFile_8 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  registerFile_9 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  registerFile_10 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  registerFile_11 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  registerFile_12 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  registerFile_13 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  registerFile_14 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  registerFile_15 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  registerFile_16 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  registerFile_17 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  registerFile_18 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  registerFile_19 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  registerFile_20 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  registerFile_21 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  registerFile_22 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  registerFile_23 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  registerFile_24 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  registerFile_25 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  registerFile_26 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  registerFile_27 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  registerFile_28 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  registerFile_29 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  registerFile_30 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  registerFile_31 = _RAND_31[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ALU(
  input  [3:0]  io_ALUCtrl,
  input  [31:0] io_A,
  input  [31:0] io_B,
  output [31:0] io_ALUOut,
  output        io_eq,
  output        io_ge,
  output        io_geu
);
  wire [4:0] shamt = io_B[4:0]; // @[ALU.scala 22:16]
  wire [31:0] _res_T_1 = $signed(io_A) & $signed(io_B); // @[ALU.scala 31:26]
  wire [31:0] _res_T_3 = $signed(io_A) | $signed(io_B); // @[ALU.scala 32:25]
  wire [31:0] _res_T_5 = $signed(io_A) ^ $signed(io_B); // @[ALU.scala 33:26]
  wire [31:0] _res_T_8 = $signed(io_A) + $signed(io_B); // @[ALU.scala 34:26]
  wire [31:0] _res_T_11 = $signed(io_A) - $signed(io_B); // @[ALU.scala 35:26]
  wire [1:0] _res_T_13 = $signed(io_A) < $signed(io_B) ? $signed(2'sh1) : $signed(2'sh0); // @[ALU.scala 36:27]
  wire [62:0] _GEN_14 = {{31{io_A[31]}},io_A}; // @[ALU.scala 37:26]
  wire [62:0] _res_T_14 = $signed(_GEN_14) << shamt; // @[ALU.scala 37:26]
  wire [1:0] _res_T_18 = io_A < io_B ? $signed(2'sh1) : $signed(2'sh0); // @[ALU.scala 38:28]
  wire [31:0] _res_T_21 = io_A >> shamt; // @[ALU.scala 39:44]
  wire [31:0] _res_T_22 = $signed(io_A) >>> shamt; // @[ALU.scala 40:26]
  wire [1:0] _res_T_27 = ~2'sh1; // @[ALU.scala 41:35]
  wire [31:0] _GEN_12 = {{30{_res_T_27[1]}},_res_T_27}; // @[ALU.scala 41:33]
  wire [31:0] _res_T_29 = $signed(_res_T_8) & $signed(_GEN_12); // @[ALU.scala 41:33]
  wire [31:0] _GEN_0 = 4'hb == io_ALUCtrl ? $signed(io_B) : $signed(32'sh0); // @[ALU.scala 30:22 24:24 42:25]
  wire [31:0] _GEN_1 = 4'ha == io_ALUCtrl ? $signed(_res_T_29) : $signed(_GEN_0); // @[ALU.scala 30:22 41:22]
  wire [31:0] _GEN_2 = 4'h9 == io_ALUCtrl ? $signed(_res_T_22) : $signed(_GEN_1); // @[ALU.scala 30:22 40:21]
  wire [31:0] _GEN_3 = 4'h8 == io_ALUCtrl ? $signed(_res_T_21) : $signed(_GEN_2); // @[ALU.scala 30:22 39:21]
  wire [31:0] _GEN_4 = 4'h7 == io_ALUCtrl ? $signed({{30{_res_T_18[1]}},_res_T_18}) : $signed(_GEN_3); // @[ALU.scala 30:22 38:22]
  wire [62:0] _GEN_5 = 4'h6 == io_ALUCtrl ? $signed(_res_T_14) : $signed({{31{_GEN_4[31]}},_GEN_4}); // @[ALU.scala 30:22 37:21]
  wire [62:0] _GEN_6 = 4'h5 == io_ALUCtrl ? $signed({{61{_res_T_13[1]}},_res_T_13}) : $signed(_GEN_5); // @[ALU.scala 30:22 36:21]
  wire [62:0] _GEN_7 = 4'h4 == io_ALUCtrl ? $signed({{31{_res_T_11[31]}},_res_T_11}) : $signed(_GEN_6); // @[ALU.scala 30:22 35:21]
  wire [62:0] _GEN_8 = 4'h3 == io_ALUCtrl ? $signed({{31{_res_T_8[31]}},_res_T_8}) : $signed(_GEN_7); // @[ALU.scala 30:22 34:21]
  wire [62:0] _GEN_9 = 4'h2 == io_ALUCtrl ? $signed({{31{_res_T_5[31]}},_res_T_5}) : $signed(_GEN_8); // @[ALU.scala 30:22 33:21]
  wire [62:0] _GEN_10 = 4'h1 == io_ALUCtrl ? $signed({{31{_res_T_3[31]}},_res_T_3}) : $signed(_GEN_9); // @[ALU.scala 30:22 32:20]
  wire [62:0] _GEN_11 = 4'h0 == io_ALUCtrl ? $signed({{31{_res_T_1[31]}},_res_T_1}) : $signed(_GEN_10); // @[ALU.scala 30:22 31:21]
  assign io_ALUOut = _GEN_11[31:0]; // @[ALU.scala 24:24]
  assign io_eq = $signed(io_A) == $signed(io_B); // @[ALU.scala 26:18]
  assign io_ge = $signed(io_A) >= $signed(io_B); // @[ALU.scala 27:18]
  assign io_geu = io_A >= io_B; // @[ALU.scala 28:26]
endmodule
module ImmGen(
  input  [31:0] io_in,
  input  [2:0]  io_format,
  output [31:0] io_out
);
  wire [11:0] _res_T_1 = io_in[31:20]; // @[ImmGen.scala 19:33]
  wire [11:0] _res_T_5 = {io_in[31:25],io_in[11:7]}; // @[ImmGen.scala 20:48]
  wire [12:0] _res_T_14 = {io_in[31],io_in[7],io_in[30:25],io_in[11:8],1'h0}; // @[ImmGen.scala 22:71]
  wire [31:0] _res_T_17 = {io_in[31:12],12'h0}; // @[ImmGen.scala 24:48]
  wire [20:0] _res_T_28 = {io_in[31],io_in[19:12],io_in[20],io_in[30:25],io_in[24:21],1'h0}; // @[ImmGen.scala 28:10]
  wire [31:0] _GEN_0 = 3'h5 == io_format ? $signed({{11{_res_T_28[20]}},_res_T_28}) : $signed(32'sh0); // @[ImmGen.scala 18:18 26:11 16:24]
  wire [31:0] _GEN_1 = 3'h4 == io_format ? $signed(_res_T_17) : $signed(_GEN_0); // @[ImmGen.scala 18:18 24:19]
  wire [31:0] _GEN_2 = 3'h3 == io_format ? $signed({{19{_res_T_14[12]}},_res_T_14}) : $signed(_GEN_1); // @[ImmGen.scala 18:18 22:11]
  wire [31:0] _GEN_3 = 3'h2 == io_format ? $signed({{20{_res_T_5[11]}},_res_T_5}) : $signed(_GEN_2); // @[ImmGen.scala 18:18 20:19]
  assign io_out = 3'h1 == io_format ? $signed({{20{_res_T_1[11]}},_res_T_1}) : $signed(_GEN_3); // @[ImmGen.scala 18:18 19:19]
endmodule
module PC(
  input         clock,
  input         reset,
  input  [31:0] io_inAddr,
  output [31:0] io_outAddr
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] io_outAddr_REG; // @[OtherComponents.scala 14:24]
  assign io_outAddr = io_outAddr_REG; // @[OtherComponents.scala 14:14]
  always @(posedge clock) begin
    if (reset) begin // @[OtherComponents.scala 14:24]
      io_outAddr_REG <= 32'h0; // @[OtherComponents.scala 14:24]
    end else begin
      io_outAddr_REG <= io_inAddr; // @[OtherComponents.scala 14:24]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  io_outAddr_REG = _RAND_0[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PCIncrementer(
  input  [31:0] io_pc,
  output [31:0] io_outAddr
);
  assign io_outAddr = io_pc + 32'h4; // @[OtherComponents.scala 23:23]
endmodule
module BranchAdder(
  input  [31:0] io_pc,
  input  [31:0] io_imm,
  output [31:0] io_outAddr
);
  assign io_outAddr = $signed(io_pc) + $signed(io_imm); // @[OtherComponents.scala 33:41]
endmodule
module PcALUMemMux(
  input         io_pcAluMem,
  input  [31:0] io_aluMem,
  input  [31:0] io_pcImm,
  output [31:0] io_out
);
  assign io_out = io_pcAluMem ? $signed(io_aluMem) : $signed(io_pcImm); // @[OtherComponents.scala 66:16]
endmodule
module Rs2ImmMux(
  input         io_rs2Imm,
  input  [31:0] io_rs2,
  input  [31:0] io_imm,
  output [31:0] io_out
);
  assign io_out = io_rs2Imm ? $signed(io_imm) : $signed(io_rs2); // @[OtherComponents.scala 44:16]
endmodule
module PcImmMux(
  input         io_pcImm,
  input  [31:0] io_pcPc4,
  input  [31:0] io_branch,
  output [31:0] io_out
);
  assign io_out = io_pcImm ? io_branch : io_pcPc4; // @[OtherComponents.scala 77:16]
endmodule
module ALUBranchMux(
  input         io_aluBranch,
  input  [31:0] io_pc4Branch,
  input  [31:0] io_ALUOut,
  output [31:0] io_out
);
  assign io_out = io_aluBranch ? io_ALUOut : io_pc4Branch; // @[OtherComponents.scala 99:16]
endmodule
module PcStallMux(
  input         io_stall,
  input  [31:0] io_next,
  input  [31:0] io_current,
  output [31:0] io_out
);
  assign io_out = io_stall ? io_next : io_current; // @[OtherComponents.scala 110:16]
endmodule
module LoadSelector(
  input  [2:0]  io_func3,
  input  [31:0] io_inData,
  output [31:0] io_outData
);
  wire [7:0] _res_T_1 = io_inData[7:0]; // @[LoadSelector.scala 19:43]
  wire [15:0] _res_T_3 = io_inData[15:0]; // @[LoadSelector.scala 20:44]
  wire [31:0] _res_T_7 = {24'h0,io_inData[7:0]}; // @[LoadSelector.scala 22:58]
  wire [31:0] _res_T_10 = {16'h0,io_inData[15:0]}; // @[LoadSelector.scala 23:59]
  wire [31:0] _GEN_0 = 3'h5 == io_func3 ? $signed(_res_T_10) : $signed(32'sh0); // @[LoadSelector.scala 18:20 16:24 23:24]
  wire [31:0] _GEN_1 = 3'h4 == io_func3 ? $signed(_res_T_7) : $signed(_GEN_0); // @[LoadSelector.scala 18:20 22:24]
  wire [31:0] _GEN_2 = 3'h2 == io_func3 ? $signed(io_inData) : $signed(_GEN_1); // @[LoadSelector.scala 18:20 21:24]
  wire [31:0] _GEN_3 = 3'h1 == io_func3 ? $signed({{16{_res_T_3[15]}},_res_T_3}) : $signed(_GEN_2); // @[LoadSelector.scala 18:20 20:24]
  assign io_outData = 3'h0 == io_func3 ? $signed({{24{_res_T_1[7]}},_res_T_1}) : $signed(_GEN_3); // @[LoadSelector.scala 18:20 19:24]
endmodule
module Core(
  input         clock,
  input         reset,
  input  [31:0] io_instr,
  input  [31:0] io_memReadData,
  input         io_valid,
  output [8:0]  io_instrAddrs,
  output [31:0] io_ALUOut,
  output [31:0] io_memWriteData,
  output        io_memRead,
  output        io_memWrite,
  output [1:0]  io_storeType
);
  wire [31:0] controlUnit_io_instr; // @[Core.scala 22:27]
  wire  controlUnit_io_eq; // @[Core.scala 22:27]
  wire  controlUnit_io_ge; // @[Core.scala 22:27]
  wire  controlUnit_io_geu; // @[Core.scala 22:27]
  wire  controlUnit_io_valid; // @[Core.scala 22:27]
  wire [2:0] controlUnit_io_format; // @[Core.scala 22:27]
  wire [3:0] controlUnit_io_ALUCtrl; // @[Core.scala 22:27]
  wire  controlUnit_io_regWrite; // @[Core.scala 22:27]
  wire  controlUnit_io_memWrite; // @[Core.scala 22:27]
  wire  controlUnit_io_memRead; // @[Core.scala 22:27]
  wire  controlUnit_io_rs2Imm; // @[Core.scala 22:27]
  wire  controlUnit_io_aluMem; // @[Core.scala 22:27]
  wire  controlUnit_io_pcAluMem; // @[Core.scala 22:27]
  wire  controlUnit_io_pcImm; // @[Core.scala 22:27]
  wire  controlUnit_io_immBranch; // @[Core.scala 22:27]
  wire  controlUnit_io_aluBranch; // @[Core.scala 22:27]
  wire  controlUnit_io_stall; // @[Core.scala 22:27]
  wire [1:0] controlUnit_io_storeType; // @[Core.scala 22:27]
  wire  registerFile_clock; // @[Core.scala 23:28]
  wire  registerFile_reset; // @[Core.scala 23:28]
  wire [4:0] registerFile_io_readAddr1; // @[Core.scala 23:28]
  wire [4:0] registerFile_io_readAddr2; // @[Core.scala 23:28]
  wire [4:0] registerFile_io_writeAddr; // @[Core.scala 23:28]
  wire [31:0] registerFile_io_writeData; // @[Core.scala 23:28]
  wire  registerFile_io_writeEn; // @[Core.scala 23:28]
  wire [31:0] registerFile_io_readData1; // @[Core.scala 23:28]
  wire [31:0] registerFile_io_readData2; // @[Core.scala 23:28]
  wire [3:0] alu_io_ALUCtrl; // @[Core.scala 24:19]
  wire [31:0] alu_io_A; // @[Core.scala 24:19]
  wire [31:0] alu_io_B; // @[Core.scala 24:19]
  wire [31:0] alu_io_ALUOut; // @[Core.scala 24:19]
  wire  alu_io_eq; // @[Core.scala 24:19]
  wire  alu_io_ge; // @[Core.scala 24:19]
  wire  alu_io_geu; // @[Core.scala 24:19]
  wire [31:0] immGen_io_in; // @[Core.scala 25:22]
  wire [2:0] immGen_io_format; // @[Core.scala 25:22]
  wire [31:0] immGen_io_out; // @[Core.scala 25:22]
  wire  pc_clock; // @[Core.scala 26:18]
  wire  pc_reset; // @[Core.scala 26:18]
  wire [31:0] pc_io_inAddr; // @[Core.scala 26:18]
  wire [31:0] pc_io_outAddr; // @[Core.scala 26:18]
  wire [31:0] pcIncrementer_io_pc; // @[Core.scala 27:29]
  wire [31:0] pcIncrementer_io_outAddr; // @[Core.scala 27:29]
  wire [31:0] branchAdder_io_pc; // @[Core.scala 28:27]
  wire [31:0] branchAdder_io_imm; // @[Core.scala 28:27]
  wire [31:0] branchAdder_io_outAddr; // @[Core.scala 28:27]
  wire  pcAluMemMux_io_pcAluMem; // @[Core.scala 29:27]
  wire [31:0] pcAluMemMux_io_aluMem; // @[Core.scala 29:27]
  wire [31:0] pcAluMemMux_io_pcImm; // @[Core.scala 29:27]
  wire [31:0] pcAluMemMux_io_out; // @[Core.scala 29:27]
  wire  rs2ImmMux_io_rs2Imm; // @[Core.scala 30:25]
  wire [31:0] rs2ImmMux_io_rs2; // @[Core.scala 30:25]
  wire [31:0] rs2ImmMux_io_imm; // @[Core.scala 30:25]
  wire [31:0] rs2ImmMux_io_out; // @[Core.scala 30:25]
  wire  pcImmMux_io_pcImm; // @[Core.scala 31:24]
  wire [31:0] pcImmMux_io_pcPc4; // @[Core.scala 31:24]
  wire [31:0] pcImmMux_io_branch; // @[Core.scala 31:24]
  wire [31:0] pcImmMux_io_out; // @[Core.scala 31:24]
  wire  aluMemMux_io_rs2Imm; // @[Core.scala 32:25]
  wire [31:0] aluMemMux_io_rs2; // @[Core.scala 32:25]
  wire [31:0] aluMemMux_io_imm; // @[Core.scala 32:25]
  wire [31:0] aluMemMux_io_out; // @[Core.scala 32:25]
  wire  immBranchMux_io_pcImm; // @[Core.scala 33:28]
  wire [31:0] immBranchMux_io_pcPc4; // @[Core.scala 33:28]
  wire [31:0] immBranchMux_io_branch; // @[Core.scala 33:28]
  wire [31:0] immBranchMux_io_out; // @[Core.scala 33:28]
  wire  aluBranchMux_io_aluBranch; // @[Core.scala 34:28]
  wire [31:0] aluBranchMux_io_pc4Branch; // @[Core.scala 34:28]
  wire [31:0] aluBranchMux_io_ALUOut; // @[Core.scala 34:28]
  wire [31:0] aluBranchMux_io_out; // @[Core.scala 34:28]
  wire  pcStall_io_stall; // @[Core.scala 35:23]
  wire [31:0] pcStall_io_next; // @[Core.scala 35:23]
  wire [31:0] pcStall_io_current; // @[Core.scala 35:23]
  wire [31:0] pcStall_io_out; // @[Core.scala 35:23]
  wire [2:0] loadSelector_io_func3; // @[Core.scala 36:28]
  wire [31:0] loadSelector_io_inData; // @[Core.scala 36:28]
  wire [31:0] loadSelector_io_outData; // @[Core.scala 36:28]
  wire [31:0] _io_instrAddrs_T = {{2'd0}, pc_io_outAddr[31:2]}; // @[Core.scala 98:35]
  ControlUnit controlUnit ( // @[Core.scala 22:27]
    .io_instr(controlUnit_io_instr),
    .io_eq(controlUnit_io_eq),
    .io_ge(controlUnit_io_ge),
    .io_geu(controlUnit_io_geu),
    .io_valid(controlUnit_io_valid),
    .io_format(controlUnit_io_format),
    .io_ALUCtrl(controlUnit_io_ALUCtrl),
    .io_regWrite(controlUnit_io_regWrite),
    .io_memWrite(controlUnit_io_memWrite),
    .io_memRead(controlUnit_io_memRead),
    .io_rs2Imm(controlUnit_io_rs2Imm),
    .io_aluMem(controlUnit_io_aluMem),
    .io_pcAluMem(controlUnit_io_pcAluMem),
    .io_pcImm(controlUnit_io_pcImm),
    .io_immBranch(controlUnit_io_immBranch),
    .io_aluBranch(controlUnit_io_aluBranch),
    .io_stall(controlUnit_io_stall),
    .io_storeType(controlUnit_io_storeType)
  );
  RegisterFile registerFile ( // @[Core.scala 23:28]
    .clock(registerFile_clock),
    .reset(registerFile_reset),
    .io_readAddr1(registerFile_io_readAddr1),
    .io_readAddr2(registerFile_io_readAddr2),
    .io_writeAddr(registerFile_io_writeAddr),
    .io_writeData(registerFile_io_writeData),
    .io_writeEn(registerFile_io_writeEn),
    .io_readData1(registerFile_io_readData1),
    .io_readData2(registerFile_io_readData2)
  );
  ALU alu ( // @[Core.scala 24:19]
    .io_ALUCtrl(alu_io_ALUCtrl),
    .io_A(alu_io_A),
    .io_B(alu_io_B),
    .io_ALUOut(alu_io_ALUOut),
    .io_eq(alu_io_eq),
    .io_ge(alu_io_ge),
    .io_geu(alu_io_geu)
  );
  ImmGen immGen ( // @[Core.scala 25:22]
    .io_in(immGen_io_in),
    .io_format(immGen_io_format),
    .io_out(immGen_io_out)
  );
  PC pc ( // @[Core.scala 26:18]
    .clock(pc_clock),
    .reset(pc_reset),
    .io_inAddr(pc_io_inAddr),
    .io_outAddr(pc_io_outAddr)
  );
  PCIncrementer pcIncrementer ( // @[Core.scala 27:29]
    .io_pc(pcIncrementer_io_pc),
    .io_outAddr(pcIncrementer_io_outAddr)
  );
  BranchAdder branchAdder ( // @[Core.scala 28:27]
    .io_pc(branchAdder_io_pc),
    .io_imm(branchAdder_io_imm),
    .io_outAddr(branchAdder_io_outAddr)
  );
  PcALUMemMux pcAluMemMux ( // @[Core.scala 29:27]
    .io_pcAluMem(pcAluMemMux_io_pcAluMem),
    .io_aluMem(pcAluMemMux_io_aluMem),
    .io_pcImm(pcAluMemMux_io_pcImm),
    .io_out(pcAluMemMux_io_out)
  );
  Rs2ImmMux rs2ImmMux ( // @[Core.scala 30:25]
    .io_rs2Imm(rs2ImmMux_io_rs2Imm),
    .io_rs2(rs2ImmMux_io_rs2),
    .io_imm(rs2ImmMux_io_imm),
    .io_out(rs2ImmMux_io_out)
  );
  PcImmMux pcImmMux ( // @[Core.scala 31:24]
    .io_pcImm(pcImmMux_io_pcImm),
    .io_pcPc4(pcImmMux_io_pcPc4),
    .io_branch(pcImmMux_io_branch),
    .io_out(pcImmMux_io_out)
  );
  Rs2ImmMux aluMemMux ( // @[Core.scala 32:25]
    .io_rs2Imm(aluMemMux_io_rs2Imm),
    .io_rs2(aluMemMux_io_rs2),
    .io_imm(aluMemMux_io_imm),
    .io_out(aluMemMux_io_out)
  );
  PcImmMux immBranchMux ( // @[Core.scala 33:28]
    .io_pcImm(immBranchMux_io_pcImm),
    .io_pcPc4(immBranchMux_io_pcPc4),
    .io_branch(immBranchMux_io_branch),
    .io_out(immBranchMux_io_out)
  );
  ALUBranchMux aluBranchMux ( // @[Core.scala 34:28]
    .io_aluBranch(aluBranchMux_io_aluBranch),
    .io_pc4Branch(aluBranchMux_io_pc4Branch),
    .io_ALUOut(aluBranchMux_io_ALUOut),
    .io_out(aluBranchMux_io_out)
  );
  PcStallMux pcStall ( // @[Core.scala 35:23]
    .io_stall(pcStall_io_stall),
    .io_next(pcStall_io_next),
    .io_current(pcStall_io_current),
    .io_out(pcStall_io_out)
  );
  LoadSelector loadSelector ( // @[Core.scala 36:28]
    .io_func3(loadSelector_io_func3),
    .io_inData(loadSelector_io_inData),
    .io_outData(loadSelector_io_outData)
  );
  assign io_instrAddrs = _io_instrAddrs_T[8:0]; // @[Core.scala 98:42]
  assign io_ALUOut = alu_io_ALUOut; // @[Core.scala 97:13]
  assign io_memWriteData = registerFile_io_readData2; // @[Core.scala 99:48]
  assign io_memRead = controlUnit_io_memRead; // @[Core.scala 95:14]
  assign io_memWrite = controlUnit_io_memWrite; // @[Core.scala 96:15]
  assign io_storeType = controlUnit_io_storeType; // @[Core.scala 100:16]
  assign controlUnit_io_instr = io_instr; // @[Core.scala 38:24]
  assign controlUnit_io_eq = alu_io_eq; // @[Core.scala 39:21]
  assign controlUnit_io_ge = alu_io_ge; // @[Core.scala 40:21]
  assign controlUnit_io_geu = alu_io_geu; // @[Core.scala 41:22]
  assign controlUnit_io_valid = io_valid; // @[Core.scala 42:24]
  assign registerFile_clock = clock;
  assign registerFile_reset = reset;
  assign registerFile_io_readAddr1 = io_instr[19:15]; // @[Core.scala 44:40]
  assign registerFile_io_readAddr2 = io_instr[24:20]; // @[Core.scala 45:40]
  assign registerFile_io_writeAddr = io_instr[11:7]; // @[Core.scala 46:40]
  assign registerFile_io_writeData = pcAluMemMux_io_out; // @[Core.scala 47:29]
  assign registerFile_io_writeEn = controlUnit_io_regWrite; // @[Core.scala 48:27]
  assign alu_io_ALUCtrl = controlUnit_io_ALUCtrl; // @[Core.scala 52:18]
  assign alu_io_A = registerFile_io_readData1; // @[Core.scala 50:12]
  assign alu_io_B = rs2ImmMux_io_out; // @[Core.scala 51:12]
  assign immGen_io_in = io_instr; // @[Core.scala 54:16]
  assign immGen_io_format = controlUnit_io_format; // @[Core.scala 55:20]
  assign pc_clock = clock;
  assign pc_reset = reset;
  assign pc_io_inAddr = pcStall_io_out; // @[Core.scala 57:16]
  assign pcIncrementer_io_pc = pc_io_outAddr; // @[Core.scala 59:23]
  assign branchAdder_io_pc = pc_io_outAddr; // @[Core.scala 61:21]
  assign branchAdder_io_imm = immGen_io_out; // @[Core.scala 62:22]
  assign pcAluMemMux_io_pcAluMem = controlUnit_io_pcAluMem; // @[Core.scala 64:27]
  assign pcAluMemMux_io_aluMem = aluMemMux_io_out; // @[Core.scala 66:25]
  assign pcAluMemMux_io_pcImm = pcImmMux_io_out; // @[Core.scala 65:24]
  assign rs2ImmMux_io_rs2Imm = controlUnit_io_rs2Imm; // @[Core.scala 68:23]
  assign rs2ImmMux_io_rs2 = registerFile_io_readData2; // @[Core.scala 70:20]
  assign rs2ImmMux_io_imm = immGen_io_out; // @[Core.scala 69:20]
  assign pcImmMux_io_pcImm = controlUnit_io_pcImm; // @[Core.scala 72:21]
  assign pcImmMux_io_pcPc4 = pcIncrementer_io_outAddr; // @[Core.scala 73:21]
  assign pcImmMux_io_branch = branchAdder_io_outAddr; // @[Core.scala 74:22]
  assign aluMemMux_io_rs2Imm = controlUnit_io_aluMem; // @[Core.scala 76:23]
  assign aluMemMux_io_rs2 = alu_io_ALUOut; // @[Core.scala 77:23]
  assign aluMemMux_io_imm = loadSelector_io_outData; // @[Core.scala 78:28]
  assign immBranchMux_io_pcImm = controlUnit_io_immBranch; // @[Core.scala 80:29]
  assign immBranchMux_io_pcPc4 = pcIncrementer_io_outAddr; // @[Core.scala 82:23]
  assign immBranchMux_io_branch = branchAdder_io_outAddr; // @[Core.scala 81:26]
  assign aluBranchMux_io_aluBranch = controlUnit_io_aluBranch; // @[Core.scala 84:29]
  assign aluBranchMux_io_pc4Branch = immBranchMux_io_out; // @[Core.scala 86:29]
  assign aluBranchMux_io_ALUOut = alu_io_ALUOut; // @[Core.scala 85:26]
  assign pcStall_io_stall = controlUnit_io_stall; // @[Core.scala 88:20]
  assign pcStall_io_next = aluBranchMux_io_out; // @[Core.scala 90:19]
  assign pcStall_io_current = pc_io_outAddr; // @[Core.scala 89:22]
  assign loadSelector_io_func3 = io_instr[14:12]; // @[Core.scala 92:36]
  assign loadSelector_io_inData = io_memReadData; // @[Core.scala 93:26]
endmodule
module L1(
  input          clock,
  input          reset,
  input  [15:0]  io_addrs,
  input  [31:0]  io_cpuWriteData,
  output [31:0]  io_cpuReadData,
  input  [1:0]   io_storeType,
  input          io_cpuWriteEn,
  output [10:0]  io_bufferAddrs,
  output [255:0] io_readBlock,
  input  [255:0] io_writeBlock,
  input          io_blockWriteEn,
  output         io_hit
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [255:0] _RAND_640;
  reg [31:0] _RAND_641;
`endif // RANDOMIZE_REG_INIT
  reg  cache_0_validBit; // @[Cache.scala 32:22]
  reg [4:0] cache_0_tag; // @[Cache.scala 32:22]
  reg [31:0] cache_0_line_0; // @[Cache.scala 32:22]
  reg [31:0] cache_0_line_1; // @[Cache.scala 32:22]
  reg [31:0] cache_0_line_2; // @[Cache.scala 32:22]
  reg [31:0] cache_0_line_3; // @[Cache.scala 32:22]
  reg [31:0] cache_0_line_4; // @[Cache.scala 32:22]
  reg [31:0] cache_0_line_5; // @[Cache.scala 32:22]
  reg [31:0] cache_0_line_6; // @[Cache.scala 32:22]
  reg [31:0] cache_0_line_7; // @[Cache.scala 32:22]
  reg  cache_1_validBit; // @[Cache.scala 32:22]
  reg [4:0] cache_1_tag; // @[Cache.scala 32:22]
  reg [31:0] cache_1_line_0; // @[Cache.scala 32:22]
  reg [31:0] cache_1_line_1; // @[Cache.scala 32:22]
  reg [31:0] cache_1_line_2; // @[Cache.scala 32:22]
  reg [31:0] cache_1_line_3; // @[Cache.scala 32:22]
  reg [31:0] cache_1_line_4; // @[Cache.scala 32:22]
  reg [31:0] cache_1_line_5; // @[Cache.scala 32:22]
  reg [31:0] cache_1_line_6; // @[Cache.scala 32:22]
  reg [31:0] cache_1_line_7; // @[Cache.scala 32:22]
  reg  cache_2_validBit; // @[Cache.scala 32:22]
  reg [4:0] cache_2_tag; // @[Cache.scala 32:22]
  reg [31:0] cache_2_line_0; // @[Cache.scala 32:22]
  reg [31:0] cache_2_line_1; // @[Cache.scala 32:22]
  reg [31:0] cache_2_line_2; // @[Cache.scala 32:22]
  reg [31:0] cache_2_line_3; // @[Cache.scala 32:22]
  reg [31:0] cache_2_line_4; // @[Cache.scala 32:22]
  reg [31:0] cache_2_line_5; // @[Cache.scala 32:22]
  reg [31:0] cache_2_line_6; // @[Cache.scala 32:22]
  reg [31:0] cache_2_line_7; // @[Cache.scala 32:22]
  reg  cache_3_validBit; // @[Cache.scala 32:22]
  reg [4:0] cache_3_tag; // @[Cache.scala 32:22]
  reg [31:0] cache_3_line_0; // @[Cache.scala 32:22]
  reg [31:0] cache_3_line_1; // @[Cache.scala 32:22]
  reg [31:0] cache_3_line_2; // @[Cache.scala 32:22]
  reg [31:0] cache_3_line_3; // @[Cache.scala 32:22]
  reg [31:0] cache_3_line_4; // @[Cache.scala 32:22]
  reg [31:0] cache_3_line_5; // @[Cache.scala 32:22]
  reg [31:0] cache_3_line_6; // @[Cache.scala 32:22]
  reg [31:0] cache_3_line_7; // @[Cache.scala 32:22]
  reg  cache_4_validBit; // @[Cache.scala 32:22]
  reg [4:0] cache_4_tag; // @[Cache.scala 32:22]
  reg [31:0] cache_4_line_0; // @[Cache.scala 32:22]
  reg [31:0] cache_4_line_1; // @[Cache.scala 32:22]
  reg [31:0] cache_4_line_2; // @[Cache.scala 32:22]
  reg [31:0] cache_4_line_3; // @[Cache.scala 32:22]
  reg [31:0] cache_4_line_4; // @[Cache.scala 32:22]
  reg [31:0] cache_4_line_5; // @[Cache.scala 32:22]
  reg [31:0] cache_4_line_6; // @[Cache.scala 32:22]
  reg [31:0] cache_4_line_7; // @[Cache.scala 32:22]
  reg  cache_5_validBit; // @[Cache.scala 32:22]
  reg [4:0] cache_5_tag; // @[Cache.scala 32:22]
  reg [31:0] cache_5_line_0; // @[Cache.scala 32:22]
  reg [31:0] cache_5_line_1; // @[Cache.scala 32:22]
  reg [31:0] cache_5_line_2; // @[Cache.scala 32:22]
  reg [31:0] cache_5_line_3; // @[Cache.scala 32:22]
  reg [31:0] cache_5_line_4; // @[Cache.scala 32:22]
  reg [31:0] cache_5_line_5; // @[Cache.scala 32:22]
  reg [31:0] cache_5_line_6; // @[Cache.scala 32:22]
  reg [31:0] cache_5_line_7; // @[Cache.scala 32:22]
  reg  cache_6_validBit; // @[Cache.scala 32:22]
  reg [4:0] cache_6_tag; // @[Cache.scala 32:22]
  reg [31:0] cache_6_line_0; // @[Cache.scala 32:22]
  reg [31:0] cache_6_line_1; // @[Cache.scala 32:22]
  reg [31:0] cache_6_line_2; // @[Cache.scala 32:22]
  reg [31:0] cache_6_line_3; // @[Cache.scala 32:22]
  reg [31:0] cache_6_line_4; // @[Cache.scala 32:22]
  reg [31:0] cache_6_line_5; // @[Cache.scala 32:22]
  reg [31:0] cache_6_line_6; // @[Cache.scala 32:22]
  reg [31:0] cache_6_line_7; // @[Cache.scala 32:22]
  reg  cache_7_validBit; // @[Cache.scala 32:22]
  reg [4:0] cache_7_tag; // @[Cache.scala 32:22]
  reg [31:0] cache_7_line_0; // @[Cache.scala 32:22]
  reg [31:0] cache_7_line_1; // @[Cache.scala 32:22]
  reg [31:0] cache_7_line_2; // @[Cache.scala 32:22]
  reg [31:0] cache_7_line_3; // @[Cache.scala 32:22]
  reg [31:0] cache_7_line_4; // @[Cache.scala 32:22]
  reg [31:0] cache_7_line_5; // @[Cache.scala 32:22]
  reg [31:0] cache_7_line_6; // @[Cache.scala 32:22]
  reg [31:0] cache_7_line_7; // @[Cache.scala 32:22]
  reg  cache_8_validBit; // @[Cache.scala 32:22]
  reg [4:0] cache_8_tag; // @[Cache.scala 32:22]
  reg [31:0] cache_8_line_0; // @[Cache.scala 32:22]
  reg [31:0] cache_8_line_1; // @[Cache.scala 32:22]
  reg [31:0] cache_8_line_2; // @[Cache.scala 32:22]
  reg [31:0] cache_8_line_3; // @[Cache.scala 32:22]
  reg [31:0] cache_8_line_4; // @[Cache.scala 32:22]
  reg [31:0] cache_8_line_5; // @[Cache.scala 32:22]
  reg [31:0] cache_8_line_6; // @[Cache.scala 32:22]
  reg [31:0] cache_8_line_7; // @[Cache.scala 32:22]
  reg  cache_9_validBit; // @[Cache.scala 32:22]
  reg [4:0] cache_9_tag; // @[Cache.scala 32:22]
  reg [31:0] cache_9_line_0; // @[Cache.scala 32:22]
  reg [31:0] cache_9_line_1; // @[Cache.scala 32:22]
  reg [31:0] cache_9_line_2; // @[Cache.scala 32:22]
  reg [31:0] cache_9_line_3; // @[Cache.scala 32:22]
  reg [31:0] cache_9_line_4; // @[Cache.scala 32:22]
  reg [31:0] cache_9_line_5; // @[Cache.scala 32:22]
  reg [31:0] cache_9_line_6; // @[Cache.scala 32:22]
  reg [31:0] cache_9_line_7; // @[Cache.scala 32:22]
  reg  cache_10_validBit; // @[Cache.scala 32:22]
  reg [4:0] cache_10_tag; // @[Cache.scala 32:22]
  reg [31:0] cache_10_line_0; // @[Cache.scala 32:22]
  reg [31:0] cache_10_line_1; // @[Cache.scala 32:22]
  reg [31:0] cache_10_line_2; // @[Cache.scala 32:22]
  reg [31:0] cache_10_line_3; // @[Cache.scala 32:22]
  reg [31:0] cache_10_line_4; // @[Cache.scala 32:22]
  reg [31:0] cache_10_line_5; // @[Cache.scala 32:22]
  reg [31:0] cache_10_line_6; // @[Cache.scala 32:22]
  reg [31:0] cache_10_line_7; // @[Cache.scala 32:22]
  reg  cache_11_validBit; // @[Cache.scala 32:22]
  reg [4:0] cache_11_tag; // @[Cache.scala 32:22]
  reg [31:0] cache_11_line_0; // @[Cache.scala 32:22]
  reg [31:0] cache_11_line_1; // @[Cache.scala 32:22]
  reg [31:0] cache_11_line_2; // @[Cache.scala 32:22]
  reg [31:0] cache_11_line_3; // @[Cache.scala 32:22]
  reg [31:0] cache_11_line_4; // @[Cache.scala 32:22]
  reg [31:0] cache_11_line_5; // @[Cache.scala 32:22]
  reg [31:0] cache_11_line_6; // @[Cache.scala 32:22]
  reg [31:0] cache_11_line_7; // @[Cache.scala 32:22]
  reg  cache_12_validBit; // @[Cache.scala 32:22]
  reg [4:0] cache_12_tag; // @[Cache.scala 32:22]
  reg [31:0] cache_12_line_0; // @[Cache.scala 32:22]
  reg [31:0] cache_12_line_1; // @[Cache.scala 32:22]
  reg [31:0] cache_12_line_2; // @[Cache.scala 32:22]
  reg [31:0] cache_12_line_3; // @[Cache.scala 32:22]
  reg [31:0] cache_12_line_4; // @[Cache.scala 32:22]
  reg [31:0] cache_12_line_5; // @[Cache.scala 32:22]
  reg [31:0] cache_12_line_6; // @[Cache.scala 32:22]
  reg [31:0] cache_12_line_7; // @[Cache.scala 32:22]
  reg  cache_13_validBit; // @[Cache.scala 32:22]
  reg [4:0] cache_13_tag; // @[Cache.scala 32:22]
  reg [31:0] cache_13_line_0; // @[Cache.scala 32:22]
  reg [31:0] cache_13_line_1; // @[Cache.scala 32:22]
  reg [31:0] cache_13_line_2; // @[Cache.scala 32:22]
  reg [31:0] cache_13_line_3; // @[Cache.scala 32:22]
  reg [31:0] cache_13_line_4; // @[Cache.scala 32:22]
  reg [31:0] cache_13_line_5; // @[Cache.scala 32:22]
  reg [31:0] cache_13_line_6; // @[Cache.scala 32:22]
  reg [31:0] cache_13_line_7; // @[Cache.scala 32:22]
  reg  cache_14_validBit; // @[Cache.scala 32:22]
  reg [4:0] cache_14_tag; // @[Cache.scala 32:22]
  reg [31:0] cache_14_line_0; // @[Cache.scala 32:22]
  reg [31:0] cache_14_line_1; // @[Cache.scala 32:22]
  reg [31:0] cache_14_line_2; // @[Cache.scala 32:22]
  reg [31:0] cache_14_line_3; // @[Cache.scala 32:22]
  reg [31:0] cache_14_line_4; // @[Cache.scala 32:22]
  reg [31:0] cache_14_line_5; // @[Cache.scala 32:22]
  reg [31:0] cache_14_line_6; // @[Cache.scala 32:22]
  reg [31:0] cache_14_line_7; // @[Cache.scala 32:22]
  reg  cache_15_validBit; // @[Cache.scala 32:22]
  reg [4:0] cache_15_tag; // @[Cache.scala 32:22]
  reg [31:0] cache_15_line_0; // @[Cache.scala 32:22]
  reg [31:0] cache_15_line_1; // @[Cache.scala 32:22]
  reg [31:0] cache_15_line_2; // @[Cache.scala 32:22]
  reg [31:0] cache_15_line_3; // @[Cache.scala 32:22]
  reg [31:0] cache_15_line_4; // @[Cache.scala 32:22]
  reg [31:0] cache_15_line_5; // @[Cache.scala 32:22]
  reg [31:0] cache_15_line_6; // @[Cache.scala 32:22]
  reg [31:0] cache_15_line_7; // @[Cache.scala 32:22]
  reg  cache_16_validBit; // @[Cache.scala 32:22]
  reg [4:0] cache_16_tag; // @[Cache.scala 32:22]
  reg [31:0] cache_16_line_0; // @[Cache.scala 32:22]
  reg [31:0] cache_16_line_1; // @[Cache.scala 32:22]
  reg [31:0] cache_16_line_2; // @[Cache.scala 32:22]
  reg [31:0] cache_16_line_3; // @[Cache.scala 32:22]
  reg [31:0] cache_16_line_4; // @[Cache.scala 32:22]
  reg [31:0] cache_16_line_5; // @[Cache.scala 32:22]
  reg [31:0] cache_16_line_6; // @[Cache.scala 32:22]
  reg [31:0] cache_16_line_7; // @[Cache.scala 32:22]
  reg  cache_17_validBit; // @[Cache.scala 32:22]
  reg [4:0] cache_17_tag; // @[Cache.scala 32:22]
  reg [31:0] cache_17_line_0; // @[Cache.scala 32:22]
  reg [31:0] cache_17_line_1; // @[Cache.scala 32:22]
  reg [31:0] cache_17_line_2; // @[Cache.scala 32:22]
  reg [31:0] cache_17_line_3; // @[Cache.scala 32:22]
  reg [31:0] cache_17_line_4; // @[Cache.scala 32:22]
  reg [31:0] cache_17_line_5; // @[Cache.scala 32:22]
  reg [31:0] cache_17_line_6; // @[Cache.scala 32:22]
  reg [31:0] cache_17_line_7; // @[Cache.scala 32:22]
  reg  cache_18_validBit; // @[Cache.scala 32:22]
  reg [4:0] cache_18_tag; // @[Cache.scala 32:22]
  reg [31:0] cache_18_line_0; // @[Cache.scala 32:22]
  reg [31:0] cache_18_line_1; // @[Cache.scala 32:22]
  reg [31:0] cache_18_line_2; // @[Cache.scala 32:22]
  reg [31:0] cache_18_line_3; // @[Cache.scala 32:22]
  reg [31:0] cache_18_line_4; // @[Cache.scala 32:22]
  reg [31:0] cache_18_line_5; // @[Cache.scala 32:22]
  reg [31:0] cache_18_line_6; // @[Cache.scala 32:22]
  reg [31:0] cache_18_line_7; // @[Cache.scala 32:22]
  reg  cache_19_validBit; // @[Cache.scala 32:22]
  reg [4:0] cache_19_tag; // @[Cache.scala 32:22]
  reg [31:0] cache_19_line_0; // @[Cache.scala 32:22]
  reg [31:0] cache_19_line_1; // @[Cache.scala 32:22]
  reg [31:0] cache_19_line_2; // @[Cache.scala 32:22]
  reg [31:0] cache_19_line_3; // @[Cache.scala 32:22]
  reg [31:0] cache_19_line_4; // @[Cache.scala 32:22]
  reg [31:0] cache_19_line_5; // @[Cache.scala 32:22]
  reg [31:0] cache_19_line_6; // @[Cache.scala 32:22]
  reg [31:0] cache_19_line_7; // @[Cache.scala 32:22]
  reg  cache_20_validBit; // @[Cache.scala 32:22]
  reg [4:0] cache_20_tag; // @[Cache.scala 32:22]
  reg [31:0] cache_20_line_0; // @[Cache.scala 32:22]
  reg [31:0] cache_20_line_1; // @[Cache.scala 32:22]
  reg [31:0] cache_20_line_2; // @[Cache.scala 32:22]
  reg [31:0] cache_20_line_3; // @[Cache.scala 32:22]
  reg [31:0] cache_20_line_4; // @[Cache.scala 32:22]
  reg [31:0] cache_20_line_5; // @[Cache.scala 32:22]
  reg [31:0] cache_20_line_6; // @[Cache.scala 32:22]
  reg [31:0] cache_20_line_7; // @[Cache.scala 32:22]
  reg  cache_21_validBit; // @[Cache.scala 32:22]
  reg [4:0] cache_21_tag; // @[Cache.scala 32:22]
  reg [31:0] cache_21_line_0; // @[Cache.scala 32:22]
  reg [31:0] cache_21_line_1; // @[Cache.scala 32:22]
  reg [31:0] cache_21_line_2; // @[Cache.scala 32:22]
  reg [31:0] cache_21_line_3; // @[Cache.scala 32:22]
  reg [31:0] cache_21_line_4; // @[Cache.scala 32:22]
  reg [31:0] cache_21_line_5; // @[Cache.scala 32:22]
  reg [31:0] cache_21_line_6; // @[Cache.scala 32:22]
  reg [31:0] cache_21_line_7; // @[Cache.scala 32:22]
  reg  cache_22_validBit; // @[Cache.scala 32:22]
  reg [4:0] cache_22_tag; // @[Cache.scala 32:22]
  reg [31:0] cache_22_line_0; // @[Cache.scala 32:22]
  reg [31:0] cache_22_line_1; // @[Cache.scala 32:22]
  reg [31:0] cache_22_line_2; // @[Cache.scala 32:22]
  reg [31:0] cache_22_line_3; // @[Cache.scala 32:22]
  reg [31:0] cache_22_line_4; // @[Cache.scala 32:22]
  reg [31:0] cache_22_line_5; // @[Cache.scala 32:22]
  reg [31:0] cache_22_line_6; // @[Cache.scala 32:22]
  reg [31:0] cache_22_line_7; // @[Cache.scala 32:22]
  reg  cache_23_validBit; // @[Cache.scala 32:22]
  reg [4:0] cache_23_tag; // @[Cache.scala 32:22]
  reg [31:0] cache_23_line_0; // @[Cache.scala 32:22]
  reg [31:0] cache_23_line_1; // @[Cache.scala 32:22]
  reg [31:0] cache_23_line_2; // @[Cache.scala 32:22]
  reg [31:0] cache_23_line_3; // @[Cache.scala 32:22]
  reg [31:0] cache_23_line_4; // @[Cache.scala 32:22]
  reg [31:0] cache_23_line_5; // @[Cache.scala 32:22]
  reg [31:0] cache_23_line_6; // @[Cache.scala 32:22]
  reg [31:0] cache_23_line_7; // @[Cache.scala 32:22]
  reg  cache_24_validBit; // @[Cache.scala 32:22]
  reg [4:0] cache_24_tag; // @[Cache.scala 32:22]
  reg [31:0] cache_24_line_0; // @[Cache.scala 32:22]
  reg [31:0] cache_24_line_1; // @[Cache.scala 32:22]
  reg [31:0] cache_24_line_2; // @[Cache.scala 32:22]
  reg [31:0] cache_24_line_3; // @[Cache.scala 32:22]
  reg [31:0] cache_24_line_4; // @[Cache.scala 32:22]
  reg [31:0] cache_24_line_5; // @[Cache.scala 32:22]
  reg [31:0] cache_24_line_6; // @[Cache.scala 32:22]
  reg [31:0] cache_24_line_7; // @[Cache.scala 32:22]
  reg  cache_25_validBit; // @[Cache.scala 32:22]
  reg [4:0] cache_25_tag; // @[Cache.scala 32:22]
  reg [31:0] cache_25_line_0; // @[Cache.scala 32:22]
  reg [31:0] cache_25_line_1; // @[Cache.scala 32:22]
  reg [31:0] cache_25_line_2; // @[Cache.scala 32:22]
  reg [31:0] cache_25_line_3; // @[Cache.scala 32:22]
  reg [31:0] cache_25_line_4; // @[Cache.scala 32:22]
  reg [31:0] cache_25_line_5; // @[Cache.scala 32:22]
  reg [31:0] cache_25_line_6; // @[Cache.scala 32:22]
  reg [31:0] cache_25_line_7; // @[Cache.scala 32:22]
  reg  cache_26_validBit; // @[Cache.scala 32:22]
  reg [4:0] cache_26_tag; // @[Cache.scala 32:22]
  reg [31:0] cache_26_line_0; // @[Cache.scala 32:22]
  reg [31:0] cache_26_line_1; // @[Cache.scala 32:22]
  reg [31:0] cache_26_line_2; // @[Cache.scala 32:22]
  reg [31:0] cache_26_line_3; // @[Cache.scala 32:22]
  reg [31:0] cache_26_line_4; // @[Cache.scala 32:22]
  reg [31:0] cache_26_line_5; // @[Cache.scala 32:22]
  reg [31:0] cache_26_line_6; // @[Cache.scala 32:22]
  reg [31:0] cache_26_line_7; // @[Cache.scala 32:22]
  reg  cache_27_validBit; // @[Cache.scala 32:22]
  reg [4:0] cache_27_tag; // @[Cache.scala 32:22]
  reg [31:0] cache_27_line_0; // @[Cache.scala 32:22]
  reg [31:0] cache_27_line_1; // @[Cache.scala 32:22]
  reg [31:0] cache_27_line_2; // @[Cache.scala 32:22]
  reg [31:0] cache_27_line_3; // @[Cache.scala 32:22]
  reg [31:0] cache_27_line_4; // @[Cache.scala 32:22]
  reg [31:0] cache_27_line_5; // @[Cache.scala 32:22]
  reg [31:0] cache_27_line_6; // @[Cache.scala 32:22]
  reg [31:0] cache_27_line_7; // @[Cache.scala 32:22]
  reg  cache_28_validBit; // @[Cache.scala 32:22]
  reg [4:0] cache_28_tag; // @[Cache.scala 32:22]
  reg [31:0] cache_28_line_0; // @[Cache.scala 32:22]
  reg [31:0] cache_28_line_1; // @[Cache.scala 32:22]
  reg [31:0] cache_28_line_2; // @[Cache.scala 32:22]
  reg [31:0] cache_28_line_3; // @[Cache.scala 32:22]
  reg [31:0] cache_28_line_4; // @[Cache.scala 32:22]
  reg [31:0] cache_28_line_5; // @[Cache.scala 32:22]
  reg [31:0] cache_28_line_6; // @[Cache.scala 32:22]
  reg [31:0] cache_28_line_7; // @[Cache.scala 32:22]
  reg  cache_29_validBit; // @[Cache.scala 32:22]
  reg [4:0] cache_29_tag; // @[Cache.scala 32:22]
  reg [31:0] cache_29_line_0; // @[Cache.scala 32:22]
  reg [31:0] cache_29_line_1; // @[Cache.scala 32:22]
  reg [31:0] cache_29_line_2; // @[Cache.scala 32:22]
  reg [31:0] cache_29_line_3; // @[Cache.scala 32:22]
  reg [31:0] cache_29_line_4; // @[Cache.scala 32:22]
  reg [31:0] cache_29_line_5; // @[Cache.scala 32:22]
  reg [31:0] cache_29_line_6; // @[Cache.scala 32:22]
  reg [31:0] cache_29_line_7; // @[Cache.scala 32:22]
  reg  cache_30_validBit; // @[Cache.scala 32:22]
  reg [4:0] cache_30_tag; // @[Cache.scala 32:22]
  reg [31:0] cache_30_line_0; // @[Cache.scala 32:22]
  reg [31:0] cache_30_line_1; // @[Cache.scala 32:22]
  reg [31:0] cache_30_line_2; // @[Cache.scala 32:22]
  reg [31:0] cache_30_line_3; // @[Cache.scala 32:22]
  reg [31:0] cache_30_line_4; // @[Cache.scala 32:22]
  reg [31:0] cache_30_line_5; // @[Cache.scala 32:22]
  reg [31:0] cache_30_line_6; // @[Cache.scala 32:22]
  reg [31:0] cache_30_line_7; // @[Cache.scala 32:22]
  reg  cache_31_validBit; // @[Cache.scala 32:22]
  reg [4:0] cache_31_tag; // @[Cache.scala 32:22]
  reg [31:0] cache_31_line_0; // @[Cache.scala 32:22]
  reg [31:0] cache_31_line_1; // @[Cache.scala 32:22]
  reg [31:0] cache_31_line_2; // @[Cache.scala 32:22]
  reg [31:0] cache_31_line_3; // @[Cache.scala 32:22]
  reg [31:0] cache_31_line_4; // @[Cache.scala 32:22]
  reg [31:0] cache_31_line_5; // @[Cache.scala 32:22]
  reg [31:0] cache_31_line_6; // @[Cache.scala 32:22]
  reg [31:0] cache_31_line_7; // @[Cache.scala 32:22]
  reg  cache_32_validBit; // @[Cache.scala 32:22]
  reg [4:0] cache_32_tag; // @[Cache.scala 32:22]
  reg [31:0] cache_32_line_0; // @[Cache.scala 32:22]
  reg [31:0] cache_32_line_1; // @[Cache.scala 32:22]
  reg [31:0] cache_32_line_2; // @[Cache.scala 32:22]
  reg [31:0] cache_32_line_3; // @[Cache.scala 32:22]
  reg [31:0] cache_32_line_4; // @[Cache.scala 32:22]
  reg [31:0] cache_32_line_5; // @[Cache.scala 32:22]
  reg [31:0] cache_32_line_6; // @[Cache.scala 32:22]
  reg [31:0] cache_32_line_7; // @[Cache.scala 32:22]
  reg  cache_33_validBit; // @[Cache.scala 32:22]
  reg [4:0] cache_33_tag; // @[Cache.scala 32:22]
  reg [31:0] cache_33_line_0; // @[Cache.scala 32:22]
  reg [31:0] cache_33_line_1; // @[Cache.scala 32:22]
  reg [31:0] cache_33_line_2; // @[Cache.scala 32:22]
  reg [31:0] cache_33_line_3; // @[Cache.scala 32:22]
  reg [31:0] cache_33_line_4; // @[Cache.scala 32:22]
  reg [31:0] cache_33_line_5; // @[Cache.scala 32:22]
  reg [31:0] cache_33_line_6; // @[Cache.scala 32:22]
  reg [31:0] cache_33_line_7; // @[Cache.scala 32:22]
  reg  cache_34_validBit; // @[Cache.scala 32:22]
  reg [4:0] cache_34_tag; // @[Cache.scala 32:22]
  reg [31:0] cache_34_line_0; // @[Cache.scala 32:22]
  reg [31:0] cache_34_line_1; // @[Cache.scala 32:22]
  reg [31:0] cache_34_line_2; // @[Cache.scala 32:22]
  reg [31:0] cache_34_line_3; // @[Cache.scala 32:22]
  reg [31:0] cache_34_line_4; // @[Cache.scala 32:22]
  reg [31:0] cache_34_line_5; // @[Cache.scala 32:22]
  reg [31:0] cache_34_line_6; // @[Cache.scala 32:22]
  reg [31:0] cache_34_line_7; // @[Cache.scala 32:22]
  reg  cache_35_validBit; // @[Cache.scala 32:22]
  reg [4:0] cache_35_tag; // @[Cache.scala 32:22]
  reg [31:0] cache_35_line_0; // @[Cache.scala 32:22]
  reg [31:0] cache_35_line_1; // @[Cache.scala 32:22]
  reg [31:0] cache_35_line_2; // @[Cache.scala 32:22]
  reg [31:0] cache_35_line_3; // @[Cache.scala 32:22]
  reg [31:0] cache_35_line_4; // @[Cache.scala 32:22]
  reg [31:0] cache_35_line_5; // @[Cache.scala 32:22]
  reg [31:0] cache_35_line_6; // @[Cache.scala 32:22]
  reg [31:0] cache_35_line_7; // @[Cache.scala 32:22]
  reg  cache_36_validBit; // @[Cache.scala 32:22]
  reg [4:0] cache_36_tag; // @[Cache.scala 32:22]
  reg [31:0] cache_36_line_0; // @[Cache.scala 32:22]
  reg [31:0] cache_36_line_1; // @[Cache.scala 32:22]
  reg [31:0] cache_36_line_2; // @[Cache.scala 32:22]
  reg [31:0] cache_36_line_3; // @[Cache.scala 32:22]
  reg [31:0] cache_36_line_4; // @[Cache.scala 32:22]
  reg [31:0] cache_36_line_5; // @[Cache.scala 32:22]
  reg [31:0] cache_36_line_6; // @[Cache.scala 32:22]
  reg [31:0] cache_36_line_7; // @[Cache.scala 32:22]
  reg  cache_37_validBit; // @[Cache.scala 32:22]
  reg [4:0] cache_37_tag; // @[Cache.scala 32:22]
  reg [31:0] cache_37_line_0; // @[Cache.scala 32:22]
  reg [31:0] cache_37_line_1; // @[Cache.scala 32:22]
  reg [31:0] cache_37_line_2; // @[Cache.scala 32:22]
  reg [31:0] cache_37_line_3; // @[Cache.scala 32:22]
  reg [31:0] cache_37_line_4; // @[Cache.scala 32:22]
  reg [31:0] cache_37_line_5; // @[Cache.scala 32:22]
  reg [31:0] cache_37_line_6; // @[Cache.scala 32:22]
  reg [31:0] cache_37_line_7; // @[Cache.scala 32:22]
  reg  cache_38_validBit; // @[Cache.scala 32:22]
  reg [4:0] cache_38_tag; // @[Cache.scala 32:22]
  reg [31:0] cache_38_line_0; // @[Cache.scala 32:22]
  reg [31:0] cache_38_line_1; // @[Cache.scala 32:22]
  reg [31:0] cache_38_line_2; // @[Cache.scala 32:22]
  reg [31:0] cache_38_line_3; // @[Cache.scala 32:22]
  reg [31:0] cache_38_line_4; // @[Cache.scala 32:22]
  reg [31:0] cache_38_line_5; // @[Cache.scala 32:22]
  reg [31:0] cache_38_line_6; // @[Cache.scala 32:22]
  reg [31:0] cache_38_line_7; // @[Cache.scala 32:22]
  reg  cache_39_validBit; // @[Cache.scala 32:22]
  reg [4:0] cache_39_tag; // @[Cache.scala 32:22]
  reg [31:0] cache_39_line_0; // @[Cache.scala 32:22]
  reg [31:0] cache_39_line_1; // @[Cache.scala 32:22]
  reg [31:0] cache_39_line_2; // @[Cache.scala 32:22]
  reg [31:0] cache_39_line_3; // @[Cache.scala 32:22]
  reg [31:0] cache_39_line_4; // @[Cache.scala 32:22]
  reg [31:0] cache_39_line_5; // @[Cache.scala 32:22]
  reg [31:0] cache_39_line_6; // @[Cache.scala 32:22]
  reg [31:0] cache_39_line_7; // @[Cache.scala 32:22]
  reg  cache_40_validBit; // @[Cache.scala 32:22]
  reg [4:0] cache_40_tag; // @[Cache.scala 32:22]
  reg [31:0] cache_40_line_0; // @[Cache.scala 32:22]
  reg [31:0] cache_40_line_1; // @[Cache.scala 32:22]
  reg [31:0] cache_40_line_2; // @[Cache.scala 32:22]
  reg [31:0] cache_40_line_3; // @[Cache.scala 32:22]
  reg [31:0] cache_40_line_4; // @[Cache.scala 32:22]
  reg [31:0] cache_40_line_5; // @[Cache.scala 32:22]
  reg [31:0] cache_40_line_6; // @[Cache.scala 32:22]
  reg [31:0] cache_40_line_7; // @[Cache.scala 32:22]
  reg  cache_41_validBit; // @[Cache.scala 32:22]
  reg [4:0] cache_41_tag; // @[Cache.scala 32:22]
  reg [31:0] cache_41_line_0; // @[Cache.scala 32:22]
  reg [31:0] cache_41_line_1; // @[Cache.scala 32:22]
  reg [31:0] cache_41_line_2; // @[Cache.scala 32:22]
  reg [31:0] cache_41_line_3; // @[Cache.scala 32:22]
  reg [31:0] cache_41_line_4; // @[Cache.scala 32:22]
  reg [31:0] cache_41_line_5; // @[Cache.scala 32:22]
  reg [31:0] cache_41_line_6; // @[Cache.scala 32:22]
  reg [31:0] cache_41_line_7; // @[Cache.scala 32:22]
  reg  cache_42_validBit; // @[Cache.scala 32:22]
  reg [4:0] cache_42_tag; // @[Cache.scala 32:22]
  reg [31:0] cache_42_line_0; // @[Cache.scala 32:22]
  reg [31:0] cache_42_line_1; // @[Cache.scala 32:22]
  reg [31:0] cache_42_line_2; // @[Cache.scala 32:22]
  reg [31:0] cache_42_line_3; // @[Cache.scala 32:22]
  reg [31:0] cache_42_line_4; // @[Cache.scala 32:22]
  reg [31:0] cache_42_line_5; // @[Cache.scala 32:22]
  reg [31:0] cache_42_line_6; // @[Cache.scala 32:22]
  reg [31:0] cache_42_line_7; // @[Cache.scala 32:22]
  reg  cache_43_validBit; // @[Cache.scala 32:22]
  reg [4:0] cache_43_tag; // @[Cache.scala 32:22]
  reg [31:0] cache_43_line_0; // @[Cache.scala 32:22]
  reg [31:0] cache_43_line_1; // @[Cache.scala 32:22]
  reg [31:0] cache_43_line_2; // @[Cache.scala 32:22]
  reg [31:0] cache_43_line_3; // @[Cache.scala 32:22]
  reg [31:0] cache_43_line_4; // @[Cache.scala 32:22]
  reg [31:0] cache_43_line_5; // @[Cache.scala 32:22]
  reg [31:0] cache_43_line_6; // @[Cache.scala 32:22]
  reg [31:0] cache_43_line_7; // @[Cache.scala 32:22]
  reg  cache_44_validBit; // @[Cache.scala 32:22]
  reg [4:0] cache_44_tag; // @[Cache.scala 32:22]
  reg [31:0] cache_44_line_0; // @[Cache.scala 32:22]
  reg [31:0] cache_44_line_1; // @[Cache.scala 32:22]
  reg [31:0] cache_44_line_2; // @[Cache.scala 32:22]
  reg [31:0] cache_44_line_3; // @[Cache.scala 32:22]
  reg [31:0] cache_44_line_4; // @[Cache.scala 32:22]
  reg [31:0] cache_44_line_5; // @[Cache.scala 32:22]
  reg [31:0] cache_44_line_6; // @[Cache.scala 32:22]
  reg [31:0] cache_44_line_7; // @[Cache.scala 32:22]
  reg  cache_45_validBit; // @[Cache.scala 32:22]
  reg [4:0] cache_45_tag; // @[Cache.scala 32:22]
  reg [31:0] cache_45_line_0; // @[Cache.scala 32:22]
  reg [31:0] cache_45_line_1; // @[Cache.scala 32:22]
  reg [31:0] cache_45_line_2; // @[Cache.scala 32:22]
  reg [31:0] cache_45_line_3; // @[Cache.scala 32:22]
  reg [31:0] cache_45_line_4; // @[Cache.scala 32:22]
  reg [31:0] cache_45_line_5; // @[Cache.scala 32:22]
  reg [31:0] cache_45_line_6; // @[Cache.scala 32:22]
  reg [31:0] cache_45_line_7; // @[Cache.scala 32:22]
  reg  cache_46_validBit; // @[Cache.scala 32:22]
  reg [4:0] cache_46_tag; // @[Cache.scala 32:22]
  reg [31:0] cache_46_line_0; // @[Cache.scala 32:22]
  reg [31:0] cache_46_line_1; // @[Cache.scala 32:22]
  reg [31:0] cache_46_line_2; // @[Cache.scala 32:22]
  reg [31:0] cache_46_line_3; // @[Cache.scala 32:22]
  reg [31:0] cache_46_line_4; // @[Cache.scala 32:22]
  reg [31:0] cache_46_line_5; // @[Cache.scala 32:22]
  reg [31:0] cache_46_line_6; // @[Cache.scala 32:22]
  reg [31:0] cache_46_line_7; // @[Cache.scala 32:22]
  reg  cache_47_validBit; // @[Cache.scala 32:22]
  reg [4:0] cache_47_tag; // @[Cache.scala 32:22]
  reg [31:0] cache_47_line_0; // @[Cache.scala 32:22]
  reg [31:0] cache_47_line_1; // @[Cache.scala 32:22]
  reg [31:0] cache_47_line_2; // @[Cache.scala 32:22]
  reg [31:0] cache_47_line_3; // @[Cache.scala 32:22]
  reg [31:0] cache_47_line_4; // @[Cache.scala 32:22]
  reg [31:0] cache_47_line_5; // @[Cache.scala 32:22]
  reg [31:0] cache_47_line_6; // @[Cache.scala 32:22]
  reg [31:0] cache_47_line_7; // @[Cache.scala 32:22]
  reg  cache_48_validBit; // @[Cache.scala 32:22]
  reg [4:0] cache_48_tag; // @[Cache.scala 32:22]
  reg [31:0] cache_48_line_0; // @[Cache.scala 32:22]
  reg [31:0] cache_48_line_1; // @[Cache.scala 32:22]
  reg [31:0] cache_48_line_2; // @[Cache.scala 32:22]
  reg [31:0] cache_48_line_3; // @[Cache.scala 32:22]
  reg [31:0] cache_48_line_4; // @[Cache.scala 32:22]
  reg [31:0] cache_48_line_5; // @[Cache.scala 32:22]
  reg [31:0] cache_48_line_6; // @[Cache.scala 32:22]
  reg [31:0] cache_48_line_7; // @[Cache.scala 32:22]
  reg  cache_49_validBit; // @[Cache.scala 32:22]
  reg [4:0] cache_49_tag; // @[Cache.scala 32:22]
  reg [31:0] cache_49_line_0; // @[Cache.scala 32:22]
  reg [31:0] cache_49_line_1; // @[Cache.scala 32:22]
  reg [31:0] cache_49_line_2; // @[Cache.scala 32:22]
  reg [31:0] cache_49_line_3; // @[Cache.scala 32:22]
  reg [31:0] cache_49_line_4; // @[Cache.scala 32:22]
  reg [31:0] cache_49_line_5; // @[Cache.scala 32:22]
  reg [31:0] cache_49_line_6; // @[Cache.scala 32:22]
  reg [31:0] cache_49_line_7; // @[Cache.scala 32:22]
  reg  cache_50_validBit; // @[Cache.scala 32:22]
  reg [4:0] cache_50_tag; // @[Cache.scala 32:22]
  reg [31:0] cache_50_line_0; // @[Cache.scala 32:22]
  reg [31:0] cache_50_line_1; // @[Cache.scala 32:22]
  reg [31:0] cache_50_line_2; // @[Cache.scala 32:22]
  reg [31:0] cache_50_line_3; // @[Cache.scala 32:22]
  reg [31:0] cache_50_line_4; // @[Cache.scala 32:22]
  reg [31:0] cache_50_line_5; // @[Cache.scala 32:22]
  reg [31:0] cache_50_line_6; // @[Cache.scala 32:22]
  reg [31:0] cache_50_line_7; // @[Cache.scala 32:22]
  reg  cache_51_validBit; // @[Cache.scala 32:22]
  reg [4:0] cache_51_tag; // @[Cache.scala 32:22]
  reg [31:0] cache_51_line_0; // @[Cache.scala 32:22]
  reg [31:0] cache_51_line_1; // @[Cache.scala 32:22]
  reg [31:0] cache_51_line_2; // @[Cache.scala 32:22]
  reg [31:0] cache_51_line_3; // @[Cache.scala 32:22]
  reg [31:0] cache_51_line_4; // @[Cache.scala 32:22]
  reg [31:0] cache_51_line_5; // @[Cache.scala 32:22]
  reg [31:0] cache_51_line_6; // @[Cache.scala 32:22]
  reg [31:0] cache_51_line_7; // @[Cache.scala 32:22]
  reg  cache_52_validBit; // @[Cache.scala 32:22]
  reg [4:0] cache_52_tag; // @[Cache.scala 32:22]
  reg [31:0] cache_52_line_0; // @[Cache.scala 32:22]
  reg [31:0] cache_52_line_1; // @[Cache.scala 32:22]
  reg [31:0] cache_52_line_2; // @[Cache.scala 32:22]
  reg [31:0] cache_52_line_3; // @[Cache.scala 32:22]
  reg [31:0] cache_52_line_4; // @[Cache.scala 32:22]
  reg [31:0] cache_52_line_5; // @[Cache.scala 32:22]
  reg [31:0] cache_52_line_6; // @[Cache.scala 32:22]
  reg [31:0] cache_52_line_7; // @[Cache.scala 32:22]
  reg  cache_53_validBit; // @[Cache.scala 32:22]
  reg [4:0] cache_53_tag; // @[Cache.scala 32:22]
  reg [31:0] cache_53_line_0; // @[Cache.scala 32:22]
  reg [31:0] cache_53_line_1; // @[Cache.scala 32:22]
  reg [31:0] cache_53_line_2; // @[Cache.scala 32:22]
  reg [31:0] cache_53_line_3; // @[Cache.scala 32:22]
  reg [31:0] cache_53_line_4; // @[Cache.scala 32:22]
  reg [31:0] cache_53_line_5; // @[Cache.scala 32:22]
  reg [31:0] cache_53_line_6; // @[Cache.scala 32:22]
  reg [31:0] cache_53_line_7; // @[Cache.scala 32:22]
  reg  cache_54_validBit; // @[Cache.scala 32:22]
  reg [4:0] cache_54_tag; // @[Cache.scala 32:22]
  reg [31:0] cache_54_line_0; // @[Cache.scala 32:22]
  reg [31:0] cache_54_line_1; // @[Cache.scala 32:22]
  reg [31:0] cache_54_line_2; // @[Cache.scala 32:22]
  reg [31:0] cache_54_line_3; // @[Cache.scala 32:22]
  reg [31:0] cache_54_line_4; // @[Cache.scala 32:22]
  reg [31:0] cache_54_line_5; // @[Cache.scala 32:22]
  reg [31:0] cache_54_line_6; // @[Cache.scala 32:22]
  reg [31:0] cache_54_line_7; // @[Cache.scala 32:22]
  reg  cache_55_validBit; // @[Cache.scala 32:22]
  reg [4:0] cache_55_tag; // @[Cache.scala 32:22]
  reg [31:0] cache_55_line_0; // @[Cache.scala 32:22]
  reg [31:0] cache_55_line_1; // @[Cache.scala 32:22]
  reg [31:0] cache_55_line_2; // @[Cache.scala 32:22]
  reg [31:0] cache_55_line_3; // @[Cache.scala 32:22]
  reg [31:0] cache_55_line_4; // @[Cache.scala 32:22]
  reg [31:0] cache_55_line_5; // @[Cache.scala 32:22]
  reg [31:0] cache_55_line_6; // @[Cache.scala 32:22]
  reg [31:0] cache_55_line_7; // @[Cache.scala 32:22]
  reg  cache_56_validBit; // @[Cache.scala 32:22]
  reg [4:0] cache_56_tag; // @[Cache.scala 32:22]
  reg [31:0] cache_56_line_0; // @[Cache.scala 32:22]
  reg [31:0] cache_56_line_1; // @[Cache.scala 32:22]
  reg [31:0] cache_56_line_2; // @[Cache.scala 32:22]
  reg [31:0] cache_56_line_3; // @[Cache.scala 32:22]
  reg [31:0] cache_56_line_4; // @[Cache.scala 32:22]
  reg [31:0] cache_56_line_5; // @[Cache.scala 32:22]
  reg [31:0] cache_56_line_6; // @[Cache.scala 32:22]
  reg [31:0] cache_56_line_7; // @[Cache.scala 32:22]
  reg  cache_57_validBit; // @[Cache.scala 32:22]
  reg [4:0] cache_57_tag; // @[Cache.scala 32:22]
  reg [31:0] cache_57_line_0; // @[Cache.scala 32:22]
  reg [31:0] cache_57_line_1; // @[Cache.scala 32:22]
  reg [31:0] cache_57_line_2; // @[Cache.scala 32:22]
  reg [31:0] cache_57_line_3; // @[Cache.scala 32:22]
  reg [31:0] cache_57_line_4; // @[Cache.scala 32:22]
  reg [31:0] cache_57_line_5; // @[Cache.scala 32:22]
  reg [31:0] cache_57_line_6; // @[Cache.scala 32:22]
  reg [31:0] cache_57_line_7; // @[Cache.scala 32:22]
  reg  cache_58_validBit; // @[Cache.scala 32:22]
  reg [4:0] cache_58_tag; // @[Cache.scala 32:22]
  reg [31:0] cache_58_line_0; // @[Cache.scala 32:22]
  reg [31:0] cache_58_line_1; // @[Cache.scala 32:22]
  reg [31:0] cache_58_line_2; // @[Cache.scala 32:22]
  reg [31:0] cache_58_line_3; // @[Cache.scala 32:22]
  reg [31:0] cache_58_line_4; // @[Cache.scala 32:22]
  reg [31:0] cache_58_line_5; // @[Cache.scala 32:22]
  reg [31:0] cache_58_line_6; // @[Cache.scala 32:22]
  reg [31:0] cache_58_line_7; // @[Cache.scala 32:22]
  reg  cache_59_validBit; // @[Cache.scala 32:22]
  reg [4:0] cache_59_tag; // @[Cache.scala 32:22]
  reg [31:0] cache_59_line_0; // @[Cache.scala 32:22]
  reg [31:0] cache_59_line_1; // @[Cache.scala 32:22]
  reg [31:0] cache_59_line_2; // @[Cache.scala 32:22]
  reg [31:0] cache_59_line_3; // @[Cache.scala 32:22]
  reg [31:0] cache_59_line_4; // @[Cache.scala 32:22]
  reg [31:0] cache_59_line_5; // @[Cache.scala 32:22]
  reg [31:0] cache_59_line_6; // @[Cache.scala 32:22]
  reg [31:0] cache_59_line_7; // @[Cache.scala 32:22]
  reg  cache_60_validBit; // @[Cache.scala 32:22]
  reg [4:0] cache_60_tag; // @[Cache.scala 32:22]
  reg [31:0] cache_60_line_0; // @[Cache.scala 32:22]
  reg [31:0] cache_60_line_1; // @[Cache.scala 32:22]
  reg [31:0] cache_60_line_2; // @[Cache.scala 32:22]
  reg [31:0] cache_60_line_3; // @[Cache.scala 32:22]
  reg [31:0] cache_60_line_4; // @[Cache.scala 32:22]
  reg [31:0] cache_60_line_5; // @[Cache.scala 32:22]
  reg [31:0] cache_60_line_6; // @[Cache.scala 32:22]
  reg [31:0] cache_60_line_7; // @[Cache.scala 32:22]
  reg  cache_61_validBit; // @[Cache.scala 32:22]
  reg [4:0] cache_61_tag; // @[Cache.scala 32:22]
  reg [31:0] cache_61_line_0; // @[Cache.scala 32:22]
  reg [31:0] cache_61_line_1; // @[Cache.scala 32:22]
  reg [31:0] cache_61_line_2; // @[Cache.scala 32:22]
  reg [31:0] cache_61_line_3; // @[Cache.scala 32:22]
  reg [31:0] cache_61_line_4; // @[Cache.scala 32:22]
  reg [31:0] cache_61_line_5; // @[Cache.scala 32:22]
  reg [31:0] cache_61_line_6; // @[Cache.scala 32:22]
  reg [31:0] cache_61_line_7; // @[Cache.scala 32:22]
  reg  cache_62_validBit; // @[Cache.scala 32:22]
  reg [4:0] cache_62_tag; // @[Cache.scala 32:22]
  reg [31:0] cache_62_line_0; // @[Cache.scala 32:22]
  reg [31:0] cache_62_line_1; // @[Cache.scala 32:22]
  reg [31:0] cache_62_line_2; // @[Cache.scala 32:22]
  reg [31:0] cache_62_line_3; // @[Cache.scala 32:22]
  reg [31:0] cache_62_line_4; // @[Cache.scala 32:22]
  reg [31:0] cache_62_line_5; // @[Cache.scala 32:22]
  reg [31:0] cache_62_line_6; // @[Cache.scala 32:22]
  reg [31:0] cache_62_line_7; // @[Cache.scala 32:22]
  reg  cache_63_validBit; // @[Cache.scala 32:22]
  reg [4:0] cache_63_tag; // @[Cache.scala 32:22]
  reg [31:0] cache_63_line_0; // @[Cache.scala 32:22]
  reg [31:0] cache_63_line_1; // @[Cache.scala 32:22]
  reg [31:0] cache_63_line_2; // @[Cache.scala 32:22]
  reg [31:0] cache_63_line_3; // @[Cache.scala 32:22]
  reg [31:0] cache_63_line_4; // @[Cache.scala 32:22]
  reg [31:0] cache_63_line_5; // @[Cache.scala 32:22]
  reg [31:0] cache_63_line_6; // @[Cache.scala 32:22]
  reg [31:0] cache_63_line_7; // @[Cache.scala 32:22]
  reg [255:0] dataBuffer; // @[Cache.scala 33:27]
  reg [15:0] addrsBuffer; // @[Cache.scala 34:28]
  wire [5:0] cacheLine = io_addrs[10:5]; // @[Cache.scala 36:27]
  wire [4:0] tag = io_addrs[15:11]; // @[Cache.scala 38:21]
  wire  _GEN_1 = 6'h1 == cacheLine ? cache_1_validBit : cache_0_validBit; // @[Cache.scala 39:{23,23}]
  wire  _GEN_2 = 6'h2 == cacheLine ? cache_2_validBit : _GEN_1; // @[Cache.scala 39:{23,23}]
  wire  _GEN_3 = 6'h3 == cacheLine ? cache_3_validBit : _GEN_2; // @[Cache.scala 39:{23,23}]
  wire  _GEN_4 = 6'h4 == cacheLine ? cache_4_validBit : _GEN_3; // @[Cache.scala 39:{23,23}]
  wire  _GEN_5 = 6'h5 == cacheLine ? cache_5_validBit : _GEN_4; // @[Cache.scala 39:{23,23}]
  wire  _GEN_6 = 6'h6 == cacheLine ? cache_6_validBit : _GEN_5; // @[Cache.scala 39:{23,23}]
  wire  _GEN_7 = 6'h7 == cacheLine ? cache_7_validBit : _GEN_6; // @[Cache.scala 39:{23,23}]
  wire  _GEN_8 = 6'h8 == cacheLine ? cache_8_validBit : _GEN_7; // @[Cache.scala 39:{23,23}]
  wire  _GEN_9 = 6'h9 == cacheLine ? cache_9_validBit : _GEN_8; // @[Cache.scala 39:{23,23}]
  wire  _GEN_10 = 6'ha == cacheLine ? cache_10_validBit : _GEN_9; // @[Cache.scala 39:{23,23}]
  wire  _GEN_11 = 6'hb == cacheLine ? cache_11_validBit : _GEN_10; // @[Cache.scala 39:{23,23}]
  wire  _GEN_12 = 6'hc == cacheLine ? cache_12_validBit : _GEN_11; // @[Cache.scala 39:{23,23}]
  wire  _GEN_13 = 6'hd == cacheLine ? cache_13_validBit : _GEN_12; // @[Cache.scala 39:{23,23}]
  wire  _GEN_14 = 6'he == cacheLine ? cache_14_validBit : _GEN_13; // @[Cache.scala 39:{23,23}]
  wire  _GEN_15 = 6'hf == cacheLine ? cache_15_validBit : _GEN_14; // @[Cache.scala 39:{23,23}]
  wire  _GEN_16 = 6'h10 == cacheLine ? cache_16_validBit : _GEN_15; // @[Cache.scala 39:{23,23}]
  wire  _GEN_17 = 6'h11 == cacheLine ? cache_17_validBit : _GEN_16; // @[Cache.scala 39:{23,23}]
  wire  _GEN_18 = 6'h12 == cacheLine ? cache_18_validBit : _GEN_17; // @[Cache.scala 39:{23,23}]
  wire  _GEN_19 = 6'h13 == cacheLine ? cache_19_validBit : _GEN_18; // @[Cache.scala 39:{23,23}]
  wire  _GEN_20 = 6'h14 == cacheLine ? cache_20_validBit : _GEN_19; // @[Cache.scala 39:{23,23}]
  wire  _GEN_21 = 6'h15 == cacheLine ? cache_21_validBit : _GEN_20; // @[Cache.scala 39:{23,23}]
  wire  _GEN_22 = 6'h16 == cacheLine ? cache_22_validBit : _GEN_21; // @[Cache.scala 39:{23,23}]
  wire  _GEN_23 = 6'h17 == cacheLine ? cache_23_validBit : _GEN_22; // @[Cache.scala 39:{23,23}]
  wire  _GEN_24 = 6'h18 == cacheLine ? cache_24_validBit : _GEN_23; // @[Cache.scala 39:{23,23}]
  wire  _GEN_25 = 6'h19 == cacheLine ? cache_25_validBit : _GEN_24; // @[Cache.scala 39:{23,23}]
  wire  _GEN_26 = 6'h1a == cacheLine ? cache_26_validBit : _GEN_25; // @[Cache.scala 39:{23,23}]
  wire  _GEN_27 = 6'h1b == cacheLine ? cache_27_validBit : _GEN_26; // @[Cache.scala 39:{23,23}]
  wire  _GEN_28 = 6'h1c == cacheLine ? cache_28_validBit : _GEN_27; // @[Cache.scala 39:{23,23}]
  wire  _GEN_29 = 6'h1d == cacheLine ? cache_29_validBit : _GEN_28; // @[Cache.scala 39:{23,23}]
  wire  _GEN_30 = 6'h1e == cacheLine ? cache_30_validBit : _GEN_29; // @[Cache.scala 39:{23,23}]
  wire  _GEN_31 = 6'h1f == cacheLine ? cache_31_validBit : _GEN_30; // @[Cache.scala 39:{23,23}]
  wire  _GEN_32 = 6'h20 == cacheLine ? cache_32_validBit : _GEN_31; // @[Cache.scala 39:{23,23}]
  wire  _GEN_33 = 6'h21 == cacheLine ? cache_33_validBit : _GEN_32; // @[Cache.scala 39:{23,23}]
  wire  _GEN_34 = 6'h22 == cacheLine ? cache_34_validBit : _GEN_33; // @[Cache.scala 39:{23,23}]
  wire  _GEN_35 = 6'h23 == cacheLine ? cache_35_validBit : _GEN_34; // @[Cache.scala 39:{23,23}]
  wire  _GEN_36 = 6'h24 == cacheLine ? cache_36_validBit : _GEN_35; // @[Cache.scala 39:{23,23}]
  wire  _GEN_37 = 6'h25 == cacheLine ? cache_37_validBit : _GEN_36; // @[Cache.scala 39:{23,23}]
  wire  _GEN_38 = 6'h26 == cacheLine ? cache_38_validBit : _GEN_37; // @[Cache.scala 39:{23,23}]
  wire  _GEN_39 = 6'h27 == cacheLine ? cache_39_validBit : _GEN_38; // @[Cache.scala 39:{23,23}]
  wire  _GEN_40 = 6'h28 == cacheLine ? cache_40_validBit : _GEN_39; // @[Cache.scala 39:{23,23}]
  wire  _GEN_41 = 6'h29 == cacheLine ? cache_41_validBit : _GEN_40; // @[Cache.scala 39:{23,23}]
  wire  _GEN_42 = 6'h2a == cacheLine ? cache_42_validBit : _GEN_41; // @[Cache.scala 39:{23,23}]
  wire  _GEN_43 = 6'h2b == cacheLine ? cache_43_validBit : _GEN_42; // @[Cache.scala 39:{23,23}]
  wire  _GEN_44 = 6'h2c == cacheLine ? cache_44_validBit : _GEN_43; // @[Cache.scala 39:{23,23}]
  wire  _GEN_45 = 6'h2d == cacheLine ? cache_45_validBit : _GEN_44; // @[Cache.scala 39:{23,23}]
  wire  _GEN_46 = 6'h2e == cacheLine ? cache_46_validBit : _GEN_45; // @[Cache.scala 39:{23,23}]
  wire  _GEN_47 = 6'h2f == cacheLine ? cache_47_validBit : _GEN_46; // @[Cache.scala 39:{23,23}]
  wire  _GEN_48 = 6'h30 == cacheLine ? cache_48_validBit : _GEN_47; // @[Cache.scala 39:{23,23}]
  wire  _GEN_49 = 6'h31 == cacheLine ? cache_49_validBit : _GEN_48; // @[Cache.scala 39:{23,23}]
  wire  _GEN_50 = 6'h32 == cacheLine ? cache_50_validBit : _GEN_49; // @[Cache.scala 39:{23,23}]
  wire  _GEN_51 = 6'h33 == cacheLine ? cache_51_validBit : _GEN_50; // @[Cache.scala 39:{23,23}]
  wire  _GEN_52 = 6'h34 == cacheLine ? cache_52_validBit : _GEN_51; // @[Cache.scala 39:{23,23}]
  wire  _GEN_53 = 6'h35 == cacheLine ? cache_53_validBit : _GEN_52; // @[Cache.scala 39:{23,23}]
  wire  _GEN_54 = 6'h36 == cacheLine ? cache_54_validBit : _GEN_53; // @[Cache.scala 39:{23,23}]
  wire  _GEN_55 = 6'h37 == cacheLine ? cache_55_validBit : _GEN_54; // @[Cache.scala 39:{23,23}]
  wire  _GEN_56 = 6'h38 == cacheLine ? cache_56_validBit : _GEN_55; // @[Cache.scala 39:{23,23}]
  wire  _GEN_57 = 6'h39 == cacheLine ? cache_57_validBit : _GEN_56; // @[Cache.scala 39:{23,23}]
  wire  _GEN_58 = 6'h3a == cacheLine ? cache_58_validBit : _GEN_57; // @[Cache.scala 39:{23,23}]
  wire  _GEN_59 = 6'h3b == cacheLine ? cache_59_validBit : _GEN_58; // @[Cache.scala 39:{23,23}]
  wire  _GEN_60 = 6'h3c == cacheLine ? cache_60_validBit : _GEN_59; // @[Cache.scala 39:{23,23}]
  wire  _GEN_61 = 6'h3d == cacheLine ? cache_61_validBit : _GEN_60; // @[Cache.scala 39:{23,23}]
  wire  _GEN_62 = 6'h3e == cacheLine ? cache_62_validBit : _GEN_61; // @[Cache.scala 39:{23,23}]
  wire  _GEN_63 = 6'h3f == cacheLine ? cache_63_validBit : _GEN_62; // @[Cache.scala 39:{23,23}]
  wire [4:0] _GEN_65 = 6'h1 == cacheLine ? cache_1_tag : cache_0_tag; // @[Cache.scala 39:{39,39}]
  wire [4:0] _GEN_66 = 6'h2 == cacheLine ? cache_2_tag : _GEN_65; // @[Cache.scala 39:{39,39}]
  wire [4:0] _GEN_67 = 6'h3 == cacheLine ? cache_3_tag : _GEN_66; // @[Cache.scala 39:{39,39}]
  wire [4:0] _GEN_68 = 6'h4 == cacheLine ? cache_4_tag : _GEN_67; // @[Cache.scala 39:{39,39}]
  wire [4:0] _GEN_69 = 6'h5 == cacheLine ? cache_5_tag : _GEN_68; // @[Cache.scala 39:{39,39}]
  wire [4:0] _GEN_70 = 6'h6 == cacheLine ? cache_6_tag : _GEN_69; // @[Cache.scala 39:{39,39}]
  wire [4:0] _GEN_71 = 6'h7 == cacheLine ? cache_7_tag : _GEN_70; // @[Cache.scala 39:{39,39}]
  wire [4:0] _GEN_72 = 6'h8 == cacheLine ? cache_8_tag : _GEN_71; // @[Cache.scala 39:{39,39}]
  wire [4:0] _GEN_73 = 6'h9 == cacheLine ? cache_9_tag : _GEN_72; // @[Cache.scala 39:{39,39}]
  wire [4:0] _GEN_74 = 6'ha == cacheLine ? cache_10_tag : _GEN_73; // @[Cache.scala 39:{39,39}]
  wire [4:0] _GEN_75 = 6'hb == cacheLine ? cache_11_tag : _GEN_74; // @[Cache.scala 39:{39,39}]
  wire [4:0] _GEN_76 = 6'hc == cacheLine ? cache_12_tag : _GEN_75; // @[Cache.scala 39:{39,39}]
  wire [4:0] _GEN_77 = 6'hd == cacheLine ? cache_13_tag : _GEN_76; // @[Cache.scala 39:{39,39}]
  wire [4:0] _GEN_78 = 6'he == cacheLine ? cache_14_tag : _GEN_77; // @[Cache.scala 39:{39,39}]
  wire [4:0] _GEN_79 = 6'hf == cacheLine ? cache_15_tag : _GEN_78; // @[Cache.scala 39:{39,39}]
  wire [4:0] _GEN_80 = 6'h10 == cacheLine ? cache_16_tag : _GEN_79; // @[Cache.scala 39:{39,39}]
  wire [4:0] _GEN_81 = 6'h11 == cacheLine ? cache_17_tag : _GEN_80; // @[Cache.scala 39:{39,39}]
  wire [4:0] _GEN_82 = 6'h12 == cacheLine ? cache_18_tag : _GEN_81; // @[Cache.scala 39:{39,39}]
  wire [4:0] _GEN_83 = 6'h13 == cacheLine ? cache_19_tag : _GEN_82; // @[Cache.scala 39:{39,39}]
  wire [4:0] _GEN_84 = 6'h14 == cacheLine ? cache_20_tag : _GEN_83; // @[Cache.scala 39:{39,39}]
  wire [4:0] _GEN_85 = 6'h15 == cacheLine ? cache_21_tag : _GEN_84; // @[Cache.scala 39:{39,39}]
  wire [4:0] _GEN_86 = 6'h16 == cacheLine ? cache_22_tag : _GEN_85; // @[Cache.scala 39:{39,39}]
  wire [4:0] _GEN_87 = 6'h17 == cacheLine ? cache_23_tag : _GEN_86; // @[Cache.scala 39:{39,39}]
  wire [4:0] _GEN_88 = 6'h18 == cacheLine ? cache_24_tag : _GEN_87; // @[Cache.scala 39:{39,39}]
  wire [4:0] _GEN_89 = 6'h19 == cacheLine ? cache_25_tag : _GEN_88; // @[Cache.scala 39:{39,39}]
  wire [4:0] _GEN_90 = 6'h1a == cacheLine ? cache_26_tag : _GEN_89; // @[Cache.scala 39:{39,39}]
  wire [4:0] _GEN_91 = 6'h1b == cacheLine ? cache_27_tag : _GEN_90; // @[Cache.scala 39:{39,39}]
  wire [4:0] _GEN_92 = 6'h1c == cacheLine ? cache_28_tag : _GEN_91; // @[Cache.scala 39:{39,39}]
  wire [4:0] _GEN_93 = 6'h1d == cacheLine ? cache_29_tag : _GEN_92; // @[Cache.scala 39:{39,39}]
  wire [4:0] _GEN_94 = 6'h1e == cacheLine ? cache_30_tag : _GEN_93; // @[Cache.scala 39:{39,39}]
  wire [4:0] _GEN_95 = 6'h1f == cacheLine ? cache_31_tag : _GEN_94; // @[Cache.scala 39:{39,39}]
  wire [4:0] _GEN_96 = 6'h20 == cacheLine ? cache_32_tag : _GEN_95; // @[Cache.scala 39:{39,39}]
  wire [4:0] _GEN_97 = 6'h21 == cacheLine ? cache_33_tag : _GEN_96; // @[Cache.scala 39:{39,39}]
  wire [4:0] _GEN_98 = 6'h22 == cacheLine ? cache_34_tag : _GEN_97; // @[Cache.scala 39:{39,39}]
  wire [4:0] _GEN_99 = 6'h23 == cacheLine ? cache_35_tag : _GEN_98; // @[Cache.scala 39:{39,39}]
  wire [4:0] _GEN_100 = 6'h24 == cacheLine ? cache_36_tag : _GEN_99; // @[Cache.scala 39:{39,39}]
  wire [4:0] _GEN_101 = 6'h25 == cacheLine ? cache_37_tag : _GEN_100; // @[Cache.scala 39:{39,39}]
  wire [4:0] _GEN_102 = 6'h26 == cacheLine ? cache_38_tag : _GEN_101; // @[Cache.scala 39:{39,39}]
  wire [4:0] _GEN_103 = 6'h27 == cacheLine ? cache_39_tag : _GEN_102; // @[Cache.scala 39:{39,39}]
  wire [4:0] _GEN_104 = 6'h28 == cacheLine ? cache_40_tag : _GEN_103; // @[Cache.scala 39:{39,39}]
  wire [4:0] _GEN_105 = 6'h29 == cacheLine ? cache_41_tag : _GEN_104; // @[Cache.scala 39:{39,39}]
  wire [4:0] _GEN_106 = 6'h2a == cacheLine ? cache_42_tag : _GEN_105; // @[Cache.scala 39:{39,39}]
  wire [4:0] _GEN_107 = 6'h2b == cacheLine ? cache_43_tag : _GEN_106; // @[Cache.scala 39:{39,39}]
  wire [4:0] _GEN_108 = 6'h2c == cacheLine ? cache_44_tag : _GEN_107; // @[Cache.scala 39:{39,39}]
  wire [4:0] _GEN_109 = 6'h2d == cacheLine ? cache_45_tag : _GEN_108; // @[Cache.scala 39:{39,39}]
  wire [4:0] _GEN_110 = 6'h2e == cacheLine ? cache_46_tag : _GEN_109; // @[Cache.scala 39:{39,39}]
  wire [4:0] _GEN_111 = 6'h2f == cacheLine ? cache_47_tag : _GEN_110; // @[Cache.scala 39:{39,39}]
  wire [4:0] _GEN_112 = 6'h30 == cacheLine ? cache_48_tag : _GEN_111; // @[Cache.scala 39:{39,39}]
  wire [4:0] _GEN_113 = 6'h31 == cacheLine ? cache_49_tag : _GEN_112; // @[Cache.scala 39:{39,39}]
  wire [4:0] _GEN_114 = 6'h32 == cacheLine ? cache_50_tag : _GEN_113; // @[Cache.scala 39:{39,39}]
  wire [4:0] _GEN_115 = 6'h33 == cacheLine ? cache_51_tag : _GEN_114; // @[Cache.scala 39:{39,39}]
  wire [4:0] _GEN_116 = 6'h34 == cacheLine ? cache_52_tag : _GEN_115; // @[Cache.scala 39:{39,39}]
  wire [4:0] _GEN_117 = 6'h35 == cacheLine ? cache_53_tag : _GEN_116; // @[Cache.scala 39:{39,39}]
  wire [4:0] _GEN_118 = 6'h36 == cacheLine ? cache_54_tag : _GEN_117; // @[Cache.scala 39:{39,39}]
  wire [4:0] _GEN_119 = 6'h37 == cacheLine ? cache_55_tag : _GEN_118; // @[Cache.scala 39:{39,39}]
  wire [4:0] _GEN_120 = 6'h38 == cacheLine ? cache_56_tag : _GEN_119; // @[Cache.scala 39:{39,39}]
  wire [4:0] _GEN_121 = 6'h39 == cacheLine ? cache_57_tag : _GEN_120; // @[Cache.scala 39:{39,39}]
  wire [4:0] _GEN_122 = 6'h3a == cacheLine ? cache_58_tag : _GEN_121; // @[Cache.scala 39:{39,39}]
  wire [4:0] _GEN_123 = 6'h3b == cacheLine ? cache_59_tag : _GEN_122; // @[Cache.scala 39:{39,39}]
  wire [4:0] _GEN_124 = 6'h3c == cacheLine ? cache_60_tag : _GEN_123; // @[Cache.scala 39:{39,39}]
  wire [4:0] _GEN_125 = 6'h3d == cacheLine ? cache_61_tag : _GEN_124; // @[Cache.scala 39:{39,39}]
  wire [4:0] _GEN_126 = 6'h3e == cacheLine ? cache_62_tag : _GEN_125; // @[Cache.scala 39:{39,39}]
  wire [4:0] _GEN_127 = 6'h3f == cacheLine ? cache_63_tag : _GEN_126; // @[Cache.scala 39:{39,39}]
  wire  hit = _GEN_63 & tag == _GEN_127; // @[Cache.scala 39:32]
  wire  _GEN_3972 = 6'h0 == cacheLine; // @[Cache.scala 40:{18,18}]
  wire  _GEN_3973 = 3'h1 == io_addrs[4:2]; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_129 = 6'h0 == cacheLine & 3'h1 == io_addrs[4:2] ? cache_0_line_1 : cache_0_line_0; // @[Cache.scala 40:{18,18}]
  wire  _GEN_3975 = 3'h2 == io_addrs[4:2]; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_130 = 6'h0 == cacheLine & 3'h2 == io_addrs[4:2] ? cache_0_line_2 : _GEN_129; // @[Cache.scala 40:{18,18}]
  wire  _GEN_3977 = 3'h3 == io_addrs[4:2]; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_131 = 6'h0 == cacheLine & 3'h3 == io_addrs[4:2] ? cache_0_line_3 : _GEN_130; // @[Cache.scala 40:{18,18}]
  wire  _GEN_3979 = 3'h4 == io_addrs[4:2]; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_132 = 6'h0 == cacheLine & 3'h4 == io_addrs[4:2] ? cache_0_line_4 : _GEN_131; // @[Cache.scala 40:{18,18}]
  wire  _GEN_3981 = 3'h5 == io_addrs[4:2]; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_133 = 6'h0 == cacheLine & 3'h5 == io_addrs[4:2] ? cache_0_line_5 : _GEN_132; // @[Cache.scala 40:{18,18}]
  wire  _GEN_3983 = 3'h6 == io_addrs[4:2]; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_134 = 6'h0 == cacheLine & 3'h6 == io_addrs[4:2] ? cache_0_line_6 : _GEN_133; // @[Cache.scala 40:{18,18}]
  wire  _GEN_3985 = 3'h7 == io_addrs[4:2]; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_135 = 6'h0 == cacheLine & 3'h7 == io_addrs[4:2] ? cache_0_line_7 : _GEN_134; // @[Cache.scala 40:{18,18}]
  wire  _GEN_3986 = 6'h1 == cacheLine; // @[Cache.scala 40:{18,18}]
  wire  _GEN_3987 = 3'h0 == io_addrs[4:2]; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_136 = 6'h1 == cacheLine & 3'h0 == io_addrs[4:2] ? cache_1_line_0 : _GEN_135; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_137 = 6'h1 == cacheLine & 3'h1 == io_addrs[4:2] ? cache_1_line_1 : _GEN_136; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_138 = 6'h1 == cacheLine & 3'h2 == io_addrs[4:2] ? cache_1_line_2 : _GEN_137; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_139 = 6'h1 == cacheLine & 3'h3 == io_addrs[4:2] ? cache_1_line_3 : _GEN_138; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_140 = 6'h1 == cacheLine & 3'h4 == io_addrs[4:2] ? cache_1_line_4 : _GEN_139; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_141 = 6'h1 == cacheLine & 3'h5 == io_addrs[4:2] ? cache_1_line_5 : _GEN_140; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_142 = 6'h1 == cacheLine & 3'h6 == io_addrs[4:2] ? cache_1_line_6 : _GEN_141; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_143 = 6'h1 == cacheLine & 3'h7 == io_addrs[4:2] ? cache_1_line_7 : _GEN_142; // @[Cache.scala 40:{18,18}]
  wire  _GEN_4002 = 6'h2 == cacheLine; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_144 = 6'h2 == cacheLine & 3'h0 == io_addrs[4:2] ? cache_2_line_0 : _GEN_143; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_145 = 6'h2 == cacheLine & 3'h1 == io_addrs[4:2] ? cache_2_line_1 : _GEN_144; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_146 = 6'h2 == cacheLine & 3'h2 == io_addrs[4:2] ? cache_2_line_2 : _GEN_145; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_147 = 6'h2 == cacheLine & 3'h3 == io_addrs[4:2] ? cache_2_line_3 : _GEN_146; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_148 = 6'h2 == cacheLine & 3'h4 == io_addrs[4:2] ? cache_2_line_4 : _GEN_147; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_149 = 6'h2 == cacheLine & 3'h5 == io_addrs[4:2] ? cache_2_line_5 : _GEN_148; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_150 = 6'h2 == cacheLine & 3'h6 == io_addrs[4:2] ? cache_2_line_6 : _GEN_149; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_151 = 6'h2 == cacheLine & 3'h7 == io_addrs[4:2] ? cache_2_line_7 : _GEN_150; // @[Cache.scala 40:{18,18}]
  wire  _GEN_4018 = 6'h3 == cacheLine; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_152 = 6'h3 == cacheLine & 3'h0 == io_addrs[4:2] ? cache_3_line_0 : _GEN_151; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_153 = 6'h3 == cacheLine & 3'h1 == io_addrs[4:2] ? cache_3_line_1 : _GEN_152; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_154 = 6'h3 == cacheLine & 3'h2 == io_addrs[4:2] ? cache_3_line_2 : _GEN_153; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_155 = 6'h3 == cacheLine & 3'h3 == io_addrs[4:2] ? cache_3_line_3 : _GEN_154; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_156 = 6'h3 == cacheLine & 3'h4 == io_addrs[4:2] ? cache_3_line_4 : _GEN_155; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_157 = 6'h3 == cacheLine & 3'h5 == io_addrs[4:2] ? cache_3_line_5 : _GEN_156; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_158 = 6'h3 == cacheLine & 3'h6 == io_addrs[4:2] ? cache_3_line_6 : _GEN_157; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_159 = 6'h3 == cacheLine & 3'h7 == io_addrs[4:2] ? cache_3_line_7 : _GEN_158; // @[Cache.scala 40:{18,18}]
  wire  _GEN_4034 = 6'h4 == cacheLine; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_160 = 6'h4 == cacheLine & 3'h0 == io_addrs[4:2] ? cache_4_line_0 : _GEN_159; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_161 = 6'h4 == cacheLine & 3'h1 == io_addrs[4:2] ? cache_4_line_1 : _GEN_160; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_162 = 6'h4 == cacheLine & 3'h2 == io_addrs[4:2] ? cache_4_line_2 : _GEN_161; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_163 = 6'h4 == cacheLine & 3'h3 == io_addrs[4:2] ? cache_4_line_3 : _GEN_162; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_164 = 6'h4 == cacheLine & 3'h4 == io_addrs[4:2] ? cache_4_line_4 : _GEN_163; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_165 = 6'h4 == cacheLine & 3'h5 == io_addrs[4:2] ? cache_4_line_5 : _GEN_164; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_166 = 6'h4 == cacheLine & 3'h6 == io_addrs[4:2] ? cache_4_line_6 : _GEN_165; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_167 = 6'h4 == cacheLine & 3'h7 == io_addrs[4:2] ? cache_4_line_7 : _GEN_166; // @[Cache.scala 40:{18,18}]
  wire  _GEN_4050 = 6'h5 == cacheLine; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_168 = 6'h5 == cacheLine & 3'h0 == io_addrs[4:2] ? cache_5_line_0 : _GEN_167; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_169 = 6'h5 == cacheLine & 3'h1 == io_addrs[4:2] ? cache_5_line_1 : _GEN_168; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_170 = 6'h5 == cacheLine & 3'h2 == io_addrs[4:2] ? cache_5_line_2 : _GEN_169; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_171 = 6'h5 == cacheLine & 3'h3 == io_addrs[4:2] ? cache_5_line_3 : _GEN_170; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_172 = 6'h5 == cacheLine & 3'h4 == io_addrs[4:2] ? cache_5_line_4 : _GEN_171; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_173 = 6'h5 == cacheLine & 3'h5 == io_addrs[4:2] ? cache_5_line_5 : _GEN_172; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_174 = 6'h5 == cacheLine & 3'h6 == io_addrs[4:2] ? cache_5_line_6 : _GEN_173; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_175 = 6'h5 == cacheLine & 3'h7 == io_addrs[4:2] ? cache_5_line_7 : _GEN_174; // @[Cache.scala 40:{18,18}]
  wire  _GEN_4066 = 6'h6 == cacheLine; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_176 = 6'h6 == cacheLine & 3'h0 == io_addrs[4:2] ? cache_6_line_0 : _GEN_175; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_177 = 6'h6 == cacheLine & 3'h1 == io_addrs[4:2] ? cache_6_line_1 : _GEN_176; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_178 = 6'h6 == cacheLine & 3'h2 == io_addrs[4:2] ? cache_6_line_2 : _GEN_177; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_179 = 6'h6 == cacheLine & 3'h3 == io_addrs[4:2] ? cache_6_line_3 : _GEN_178; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_180 = 6'h6 == cacheLine & 3'h4 == io_addrs[4:2] ? cache_6_line_4 : _GEN_179; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_181 = 6'h6 == cacheLine & 3'h5 == io_addrs[4:2] ? cache_6_line_5 : _GEN_180; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_182 = 6'h6 == cacheLine & 3'h6 == io_addrs[4:2] ? cache_6_line_6 : _GEN_181; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_183 = 6'h6 == cacheLine & 3'h7 == io_addrs[4:2] ? cache_6_line_7 : _GEN_182; // @[Cache.scala 40:{18,18}]
  wire  _GEN_4082 = 6'h7 == cacheLine; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_184 = 6'h7 == cacheLine & 3'h0 == io_addrs[4:2] ? cache_7_line_0 : _GEN_183; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_185 = 6'h7 == cacheLine & 3'h1 == io_addrs[4:2] ? cache_7_line_1 : _GEN_184; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_186 = 6'h7 == cacheLine & 3'h2 == io_addrs[4:2] ? cache_7_line_2 : _GEN_185; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_187 = 6'h7 == cacheLine & 3'h3 == io_addrs[4:2] ? cache_7_line_3 : _GEN_186; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_188 = 6'h7 == cacheLine & 3'h4 == io_addrs[4:2] ? cache_7_line_4 : _GEN_187; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_189 = 6'h7 == cacheLine & 3'h5 == io_addrs[4:2] ? cache_7_line_5 : _GEN_188; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_190 = 6'h7 == cacheLine & 3'h6 == io_addrs[4:2] ? cache_7_line_6 : _GEN_189; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_191 = 6'h7 == cacheLine & 3'h7 == io_addrs[4:2] ? cache_7_line_7 : _GEN_190; // @[Cache.scala 40:{18,18}]
  wire  _GEN_4098 = 6'h8 == cacheLine; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_192 = 6'h8 == cacheLine & 3'h0 == io_addrs[4:2] ? cache_8_line_0 : _GEN_191; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_193 = 6'h8 == cacheLine & 3'h1 == io_addrs[4:2] ? cache_8_line_1 : _GEN_192; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_194 = 6'h8 == cacheLine & 3'h2 == io_addrs[4:2] ? cache_8_line_2 : _GEN_193; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_195 = 6'h8 == cacheLine & 3'h3 == io_addrs[4:2] ? cache_8_line_3 : _GEN_194; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_196 = 6'h8 == cacheLine & 3'h4 == io_addrs[4:2] ? cache_8_line_4 : _GEN_195; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_197 = 6'h8 == cacheLine & 3'h5 == io_addrs[4:2] ? cache_8_line_5 : _GEN_196; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_198 = 6'h8 == cacheLine & 3'h6 == io_addrs[4:2] ? cache_8_line_6 : _GEN_197; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_199 = 6'h8 == cacheLine & 3'h7 == io_addrs[4:2] ? cache_8_line_7 : _GEN_198; // @[Cache.scala 40:{18,18}]
  wire  _GEN_4114 = 6'h9 == cacheLine; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_200 = 6'h9 == cacheLine & 3'h0 == io_addrs[4:2] ? cache_9_line_0 : _GEN_199; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_201 = 6'h9 == cacheLine & 3'h1 == io_addrs[4:2] ? cache_9_line_1 : _GEN_200; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_202 = 6'h9 == cacheLine & 3'h2 == io_addrs[4:2] ? cache_9_line_2 : _GEN_201; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_203 = 6'h9 == cacheLine & 3'h3 == io_addrs[4:2] ? cache_9_line_3 : _GEN_202; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_204 = 6'h9 == cacheLine & 3'h4 == io_addrs[4:2] ? cache_9_line_4 : _GEN_203; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_205 = 6'h9 == cacheLine & 3'h5 == io_addrs[4:2] ? cache_9_line_5 : _GEN_204; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_206 = 6'h9 == cacheLine & 3'h6 == io_addrs[4:2] ? cache_9_line_6 : _GEN_205; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_207 = 6'h9 == cacheLine & 3'h7 == io_addrs[4:2] ? cache_9_line_7 : _GEN_206; // @[Cache.scala 40:{18,18}]
  wire  _GEN_4130 = 6'ha == cacheLine; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_208 = 6'ha == cacheLine & 3'h0 == io_addrs[4:2] ? cache_10_line_0 : _GEN_207; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_209 = 6'ha == cacheLine & 3'h1 == io_addrs[4:2] ? cache_10_line_1 : _GEN_208; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_210 = 6'ha == cacheLine & 3'h2 == io_addrs[4:2] ? cache_10_line_2 : _GEN_209; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_211 = 6'ha == cacheLine & 3'h3 == io_addrs[4:2] ? cache_10_line_3 : _GEN_210; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_212 = 6'ha == cacheLine & 3'h4 == io_addrs[4:2] ? cache_10_line_4 : _GEN_211; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_213 = 6'ha == cacheLine & 3'h5 == io_addrs[4:2] ? cache_10_line_5 : _GEN_212; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_214 = 6'ha == cacheLine & 3'h6 == io_addrs[4:2] ? cache_10_line_6 : _GEN_213; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_215 = 6'ha == cacheLine & 3'h7 == io_addrs[4:2] ? cache_10_line_7 : _GEN_214; // @[Cache.scala 40:{18,18}]
  wire  _GEN_4146 = 6'hb == cacheLine; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_216 = 6'hb == cacheLine & 3'h0 == io_addrs[4:2] ? cache_11_line_0 : _GEN_215; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_217 = 6'hb == cacheLine & 3'h1 == io_addrs[4:2] ? cache_11_line_1 : _GEN_216; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_218 = 6'hb == cacheLine & 3'h2 == io_addrs[4:2] ? cache_11_line_2 : _GEN_217; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_219 = 6'hb == cacheLine & 3'h3 == io_addrs[4:2] ? cache_11_line_3 : _GEN_218; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_220 = 6'hb == cacheLine & 3'h4 == io_addrs[4:2] ? cache_11_line_4 : _GEN_219; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_221 = 6'hb == cacheLine & 3'h5 == io_addrs[4:2] ? cache_11_line_5 : _GEN_220; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_222 = 6'hb == cacheLine & 3'h6 == io_addrs[4:2] ? cache_11_line_6 : _GEN_221; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_223 = 6'hb == cacheLine & 3'h7 == io_addrs[4:2] ? cache_11_line_7 : _GEN_222; // @[Cache.scala 40:{18,18}]
  wire  _GEN_4162 = 6'hc == cacheLine; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_224 = 6'hc == cacheLine & 3'h0 == io_addrs[4:2] ? cache_12_line_0 : _GEN_223; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_225 = 6'hc == cacheLine & 3'h1 == io_addrs[4:2] ? cache_12_line_1 : _GEN_224; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_226 = 6'hc == cacheLine & 3'h2 == io_addrs[4:2] ? cache_12_line_2 : _GEN_225; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_227 = 6'hc == cacheLine & 3'h3 == io_addrs[4:2] ? cache_12_line_3 : _GEN_226; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_228 = 6'hc == cacheLine & 3'h4 == io_addrs[4:2] ? cache_12_line_4 : _GEN_227; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_229 = 6'hc == cacheLine & 3'h5 == io_addrs[4:2] ? cache_12_line_5 : _GEN_228; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_230 = 6'hc == cacheLine & 3'h6 == io_addrs[4:2] ? cache_12_line_6 : _GEN_229; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_231 = 6'hc == cacheLine & 3'h7 == io_addrs[4:2] ? cache_12_line_7 : _GEN_230; // @[Cache.scala 40:{18,18}]
  wire  _GEN_4178 = 6'hd == cacheLine; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_232 = 6'hd == cacheLine & 3'h0 == io_addrs[4:2] ? cache_13_line_0 : _GEN_231; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_233 = 6'hd == cacheLine & 3'h1 == io_addrs[4:2] ? cache_13_line_1 : _GEN_232; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_234 = 6'hd == cacheLine & 3'h2 == io_addrs[4:2] ? cache_13_line_2 : _GEN_233; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_235 = 6'hd == cacheLine & 3'h3 == io_addrs[4:2] ? cache_13_line_3 : _GEN_234; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_236 = 6'hd == cacheLine & 3'h4 == io_addrs[4:2] ? cache_13_line_4 : _GEN_235; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_237 = 6'hd == cacheLine & 3'h5 == io_addrs[4:2] ? cache_13_line_5 : _GEN_236; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_238 = 6'hd == cacheLine & 3'h6 == io_addrs[4:2] ? cache_13_line_6 : _GEN_237; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_239 = 6'hd == cacheLine & 3'h7 == io_addrs[4:2] ? cache_13_line_7 : _GEN_238; // @[Cache.scala 40:{18,18}]
  wire  _GEN_4194 = 6'he == cacheLine; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_240 = 6'he == cacheLine & 3'h0 == io_addrs[4:2] ? cache_14_line_0 : _GEN_239; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_241 = 6'he == cacheLine & 3'h1 == io_addrs[4:2] ? cache_14_line_1 : _GEN_240; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_242 = 6'he == cacheLine & 3'h2 == io_addrs[4:2] ? cache_14_line_2 : _GEN_241; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_243 = 6'he == cacheLine & 3'h3 == io_addrs[4:2] ? cache_14_line_3 : _GEN_242; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_244 = 6'he == cacheLine & 3'h4 == io_addrs[4:2] ? cache_14_line_4 : _GEN_243; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_245 = 6'he == cacheLine & 3'h5 == io_addrs[4:2] ? cache_14_line_5 : _GEN_244; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_246 = 6'he == cacheLine & 3'h6 == io_addrs[4:2] ? cache_14_line_6 : _GEN_245; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_247 = 6'he == cacheLine & 3'h7 == io_addrs[4:2] ? cache_14_line_7 : _GEN_246; // @[Cache.scala 40:{18,18}]
  wire  _GEN_4210 = 6'hf == cacheLine; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_248 = 6'hf == cacheLine & 3'h0 == io_addrs[4:2] ? cache_15_line_0 : _GEN_247; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_249 = 6'hf == cacheLine & 3'h1 == io_addrs[4:2] ? cache_15_line_1 : _GEN_248; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_250 = 6'hf == cacheLine & 3'h2 == io_addrs[4:2] ? cache_15_line_2 : _GEN_249; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_251 = 6'hf == cacheLine & 3'h3 == io_addrs[4:2] ? cache_15_line_3 : _GEN_250; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_252 = 6'hf == cacheLine & 3'h4 == io_addrs[4:2] ? cache_15_line_4 : _GEN_251; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_253 = 6'hf == cacheLine & 3'h5 == io_addrs[4:2] ? cache_15_line_5 : _GEN_252; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_254 = 6'hf == cacheLine & 3'h6 == io_addrs[4:2] ? cache_15_line_6 : _GEN_253; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_255 = 6'hf == cacheLine & 3'h7 == io_addrs[4:2] ? cache_15_line_7 : _GEN_254; // @[Cache.scala 40:{18,18}]
  wire  _GEN_4226 = 6'h10 == cacheLine; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_256 = 6'h10 == cacheLine & 3'h0 == io_addrs[4:2] ? cache_16_line_0 : _GEN_255; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_257 = 6'h10 == cacheLine & 3'h1 == io_addrs[4:2] ? cache_16_line_1 : _GEN_256; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_258 = 6'h10 == cacheLine & 3'h2 == io_addrs[4:2] ? cache_16_line_2 : _GEN_257; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_259 = 6'h10 == cacheLine & 3'h3 == io_addrs[4:2] ? cache_16_line_3 : _GEN_258; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_260 = 6'h10 == cacheLine & 3'h4 == io_addrs[4:2] ? cache_16_line_4 : _GEN_259; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_261 = 6'h10 == cacheLine & 3'h5 == io_addrs[4:2] ? cache_16_line_5 : _GEN_260; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_262 = 6'h10 == cacheLine & 3'h6 == io_addrs[4:2] ? cache_16_line_6 : _GEN_261; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_263 = 6'h10 == cacheLine & 3'h7 == io_addrs[4:2] ? cache_16_line_7 : _GEN_262; // @[Cache.scala 40:{18,18}]
  wire  _GEN_4242 = 6'h11 == cacheLine; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_264 = 6'h11 == cacheLine & 3'h0 == io_addrs[4:2] ? cache_17_line_0 : _GEN_263; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_265 = 6'h11 == cacheLine & 3'h1 == io_addrs[4:2] ? cache_17_line_1 : _GEN_264; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_266 = 6'h11 == cacheLine & 3'h2 == io_addrs[4:2] ? cache_17_line_2 : _GEN_265; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_267 = 6'h11 == cacheLine & 3'h3 == io_addrs[4:2] ? cache_17_line_3 : _GEN_266; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_268 = 6'h11 == cacheLine & 3'h4 == io_addrs[4:2] ? cache_17_line_4 : _GEN_267; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_269 = 6'h11 == cacheLine & 3'h5 == io_addrs[4:2] ? cache_17_line_5 : _GEN_268; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_270 = 6'h11 == cacheLine & 3'h6 == io_addrs[4:2] ? cache_17_line_6 : _GEN_269; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_271 = 6'h11 == cacheLine & 3'h7 == io_addrs[4:2] ? cache_17_line_7 : _GEN_270; // @[Cache.scala 40:{18,18}]
  wire  _GEN_4258 = 6'h12 == cacheLine; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_272 = 6'h12 == cacheLine & 3'h0 == io_addrs[4:2] ? cache_18_line_0 : _GEN_271; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_273 = 6'h12 == cacheLine & 3'h1 == io_addrs[4:2] ? cache_18_line_1 : _GEN_272; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_274 = 6'h12 == cacheLine & 3'h2 == io_addrs[4:2] ? cache_18_line_2 : _GEN_273; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_275 = 6'h12 == cacheLine & 3'h3 == io_addrs[4:2] ? cache_18_line_3 : _GEN_274; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_276 = 6'h12 == cacheLine & 3'h4 == io_addrs[4:2] ? cache_18_line_4 : _GEN_275; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_277 = 6'h12 == cacheLine & 3'h5 == io_addrs[4:2] ? cache_18_line_5 : _GEN_276; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_278 = 6'h12 == cacheLine & 3'h6 == io_addrs[4:2] ? cache_18_line_6 : _GEN_277; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_279 = 6'h12 == cacheLine & 3'h7 == io_addrs[4:2] ? cache_18_line_7 : _GEN_278; // @[Cache.scala 40:{18,18}]
  wire  _GEN_4274 = 6'h13 == cacheLine; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_280 = 6'h13 == cacheLine & 3'h0 == io_addrs[4:2] ? cache_19_line_0 : _GEN_279; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_281 = 6'h13 == cacheLine & 3'h1 == io_addrs[4:2] ? cache_19_line_1 : _GEN_280; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_282 = 6'h13 == cacheLine & 3'h2 == io_addrs[4:2] ? cache_19_line_2 : _GEN_281; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_283 = 6'h13 == cacheLine & 3'h3 == io_addrs[4:2] ? cache_19_line_3 : _GEN_282; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_284 = 6'h13 == cacheLine & 3'h4 == io_addrs[4:2] ? cache_19_line_4 : _GEN_283; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_285 = 6'h13 == cacheLine & 3'h5 == io_addrs[4:2] ? cache_19_line_5 : _GEN_284; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_286 = 6'h13 == cacheLine & 3'h6 == io_addrs[4:2] ? cache_19_line_6 : _GEN_285; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_287 = 6'h13 == cacheLine & 3'h7 == io_addrs[4:2] ? cache_19_line_7 : _GEN_286; // @[Cache.scala 40:{18,18}]
  wire  _GEN_4290 = 6'h14 == cacheLine; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_288 = 6'h14 == cacheLine & 3'h0 == io_addrs[4:2] ? cache_20_line_0 : _GEN_287; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_289 = 6'h14 == cacheLine & 3'h1 == io_addrs[4:2] ? cache_20_line_1 : _GEN_288; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_290 = 6'h14 == cacheLine & 3'h2 == io_addrs[4:2] ? cache_20_line_2 : _GEN_289; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_291 = 6'h14 == cacheLine & 3'h3 == io_addrs[4:2] ? cache_20_line_3 : _GEN_290; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_292 = 6'h14 == cacheLine & 3'h4 == io_addrs[4:2] ? cache_20_line_4 : _GEN_291; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_293 = 6'h14 == cacheLine & 3'h5 == io_addrs[4:2] ? cache_20_line_5 : _GEN_292; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_294 = 6'h14 == cacheLine & 3'h6 == io_addrs[4:2] ? cache_20_line_6 : _GEN_293; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_295 = 6'h14 == cacheLine & 3'h7 == io_addrs[4:2] ? cache_20_line_7 : _GEN_294; // @[Cache.scala 40:{18,18}]
  wire  _GEN_4306 = 6'h15 == cacheLine; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_296 = 6'h15 == cacheLine & 3'h0 == io_addrs[4:2] ? cache_21_line_0 : _GEN_295; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_297 = 6'h15 == cacheLine & 3'h1 == io_addrs[4:2] ? cache_21_line_1 : _GEN_296; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_298 = 6'h15 == cacheLine & 3'h2 == io_addrs[4:2] ? cache_21_line_2 : _GEN_297; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_299 = 6'h15 == cacheLine & 3'h3 == io_addrs[4:2] ? cache_21_line_3 : _GEN_298; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_300 = 6'h15 == cacheLine & 3'h4 == io_addrs[4:2] ? cache_21_line_4 : _GEN_299; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_301 = 6'h15 == cacheLine & 3'h5 == io_addrs[4:2] ? cache_21_line_5 : _GEN_300; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_302 = 6'h15 == cacheLine & 3'h6 == io_addrs[4:2] ? cache_21_line_6 : _GEN_301; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_303 = 6'h15 == cacheLine & 3'h7 == io_addrs[4:2] ? cache_21_line_7 : _GEN_302; // @[Cache.scala 40:{18,18}]
  wire  _GEN_4322 = 6'h16 == cacheLine; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_304 = 6'h16 == cacheLine & 3'h0 == io_addrs[4:2] ? cache_22_line_0 : _GEN_303; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_305 = 6'h16 == cacheLine & 3'h1 == io_addrs[4:2] ? cache_22_line_1 : _GEN_304; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_306 = 6'h16 == cacheLine & 3'h2 == io_addrs[4:2] ? cache_22_line_2 : _GEN_305; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_307 = 6'h16 == cacheLine & 3'h3 == io_addrs[4:2] ? cache_22_line_3 : _GEN_306; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_308 = 6'h16 == cacheLine & 3'h4 == io_addrs[4:2] ? cache_22_line_4 : _GEN_307; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_309 = 6'h16 == cacheLine & 3'h5 == io_addrs[4:2] ? cache_22_line_5 : _GEN_308; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_310 = 6'h16 == cacheLine & 3'h6 == io_addrs[4:2] ? cache_22_line_6 : _GEN_309; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_311 = 6'h16 == cacheLine & 3'h7 == io_addrs[4:2] ? cache_22_line_7 : _GEN_310; // @[Cache.scala 40:{18,18}]
  wire  _GEN_4338 = 6'h17 == cacheLine; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_312 = 6'h17 == cacheLine & 3'h0 == io_addrs[4:2] ? cache_23_line_0 : _GEN_311; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_313 = 6'h17 == cacheLine & 3'h1 == io_addrs[4:2] ? cache_23_line_1 : _GEN_312; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_314 = 6'h17 == cacheLine & 3'h2 == io_addrs[4:2] ? cache_23_line_2 : _GEN_313; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_315 = 6'h17 == cacheLine & 3'h3 == io_addrs[4:2] ? cache_23_line_3 : _GEN_314; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_316 = 6'h17 == cacheLine & 3'h4 == io_addrs[4:2] ? cache_23_line_4 : _GEN_315; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_317 = 6'h17 == cacheLine & 3'h5 == io_addrs[4:2] ? cache_23_line_5 : _GEN_316; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_318 = 6'h17 == cacheLine & 3'h6 == io_addrs[4:2] ? cache_23_line_6 : _GEN_317; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_319 = 6'h17 == cacheLine & 3'h7 == io_addrs[4:2] ? cache_23_line_7 : _GEN_318; // @[Cache.scala 40:{18,18}]
  wire  _GEN_4354 = 6'h18 == cacheLine; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_320 = 6'h18 == cacheLine & 3'h0 == io_addrs[4:2] ? cache_24_line_0 : _GEN_319; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_321 = 6'h18 == cacheLine & 3'h1 == io_addrs[4:2] ? cache_24_line_1 : _GEN_320; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_322 = 6'h18 == cacheLine & 3'h2 == io_addrs[4:2] ? cache_24_line_2 : _GEN_321; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_323 = 6'h18 == cacheLine & 3'h3 == io_addrs[4:2] ? cache_24_line_3 : _GEN_322; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_324 = 6'h18 == cacheLine & 3'h4 == io_addrs[4:2] ? cache_24_line_4 : _GEN_323; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_325 = 6'h18 == cacheLine & 3'h5 == io_addrs[4:2] ? cache_24_line_5 : _GEN_324; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_326 = 6'h18 == cacheLine & 3'h6 == io_addrs[4:2] ? cache_24_line_6 : _GEN_325; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_327 = 6'h18 == cacheLine & 3'h7 == io_addrs[4:2] ? cache_24_line_7 : _GEN_326; // @[Cache.scala 40:{18,18}]
  wire  _GEN_4370 = 6'h19 == cacheLine; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_328 = 6'h19 == cacheLine & 3'h0 == io_addrs[4:2] ? cache_25_line_0 : _GEN_327; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_329 = 6'h19 == cacheLine & 3'h1 == io_addrs[4:2] ? cache_25_line_1 : _GEN_328; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_330 = 6'h19 == cacheLine & 3'h2 == io_addrs[4:2] ? cache_25_line_2 : _GEN_329; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_331 = 6'h19 == cacheLine & 3'h3 == io_addrs[4:2] ? cache_25_line_3 : _GEN_330; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_332 = 6'h19 == cacheLine & 3'h4 == io_addrs[4:2] ? cache_25_line_4 : _GEN_331; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_333 = 6'h19 == cacheLine & 3'h5 == io_addrs[4:2] ? cache_25_line_5 : _GEN_332; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_334 = 6'h19 == cacheLine & 3'h6 == io_addrs[4:2] ? cache_25_line_6 : _GEN_333; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_335 = 6'h19 == cacheLine & 3'h7 == io_addrs[4:2] ? cache_25_line_7 : _GEN_334; // @[Cache.scala 40:{18,18}]
  wire  _GEN_4386 = 6'h1a == cacheLine; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_336 = 6'h1a == cacheLine & 3'h0 == io_addrs[4:2] ? cache_26_line_0 : _GEN_335; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_337 = 6'h1a == cacheLine & 3'h1 == io_addrs[4:2] ? cache_26_line_1 : _GEN_336; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_338 = 6'h1a == cacheLine & 3'h2 == io_addrs[4:2] ? cache_26_line_2 : _GEN_337; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_339 = 6'h1a == cacheLine & 3'h3 == io_addrs[4:2] ? cache_26_line_3 : _GEN_338; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_340 = 6'h1a == cacheLine & 3'h4 == io_addrs[4:2] ? cache_26_line_4 : _GEN_339; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_341 = 6'h1a == cacheLine & 3'h5 == io_addrs[4:2] ? cache_26_line_5 : _GEN_340; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_342 = 6'h1a == cacheLine & 3'h6 == io_addrs[4:2] ? cache_26_line_6 : _GEN_341; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_343 = 6'h1a == cacheLine & 3'h7 == io_addrs[4:2] ? cache_26_line_7 : _GEN_342; // @[Cache.scala 40:{18,18}]
  wire  _GEN_4402 = 6'h1b == cacheLine; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_344 = 6'h1b == cacheLine & 3'h0 == io_addrs[4:2] ? cache_27_line_0 : _GEN_343; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_345 = 6'h1b == cacheLine & 3'h1 == io_addrs[4:2] ? cache_27_line_1 : _GEN_344; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_346 = 6'h1b == cacheLine & 3'h2 == io_addrs[4:2] ? cache_27_line_2 : _GEN_345; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_347 = 6'h1b == cacheLine & 3'h3 == io_addrs[4:2] ? cache_27_line_3 : _GEN_346; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_348 = 6'h1b == cacheLine & 3'h4 == io_addrs[4:2] ? cache_27_line_4 : _GEN_347; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_349 = 6'h1b == cacheLine & 3'h5 == io_addrs[4:2] ? cache_27_line_5 : _GEN_348; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_350 = 6'h1b == cacheLine & 3'h6 == io_addrs[4:2] ? cache_27_line_6 : _GEN_349; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_351 = 6'h1b == cacheLine & 3'h7 == io_addrs[4:2] ? cache_27_line_7 : _GEN_350; // @[Cache.scala 40:{18,18}]
  wire  _GEN_4418 = 6'h1c == cacheLine; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_352 = 6'h1c == cacheLine & 3'h0 == io_addrs[4:2] ? cache_28_line_0 : _GEN_351; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_353 = 6'h1c == cacheLine & 3'h1 == io_addrs[4:2] ? cache_28_line_1 : _GEN_352; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_354 = 6'h1c == cacheLine & 3'h2 == io_addrs[4:2] ? cache_28_line_2 : _GEN_353; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_355 = 6'h1c == cacheLine & 3'h3 == io_addrs[4:2] ? cache_28_line_3 : _GEN_354; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_356 = 6'h1c == cacheLine & 3'h4 == io_addrs[4:2] ? cache_28_line_4 : _GEN_355; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_357 = 6'h1c == cacheLine & 3'h5 == io_addrs[4:2] ? cache_28_line_5 : _GEN_356; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_358 = 6'h1c == cacheLine & 3'h6 == io_addrs[4:2] ? cache_28_line_6 : _GEN_357; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_359 = 6'h1c == cacheLine & 3'h7 == io_addrs[4:2] ? cache_28_line_7 : _GEN_358; // @[Cache.scala 40:{18,18}]
  wire  _GEN_4434 = 6'h1d == cacheLine; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_360 = 6'h1d == cacheLine & 3'h0 == io_addrs[4:2] ? cache_29_line_0 : _GEN_359; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_361 = 6'h1d == cacheLine & 3'h1 == io_addrs[4:2] ? cache_29_line_1 : _GEN_360; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_362 = 6'h1d == cacheLine & 3'h2 == io_addrs[4:2] ? cache_29_line_2 : _GEN_361; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_363 = 6'h1d == cacheLine & 3'h3 == io_addrs[4:2] ? cache_29_line_3 : _GEN_362; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_364 = 6'h1d == cacheLine & 3'h4 == io_addrs[4:2] ? cache_29_line_4 : _GEN_363; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_365 = 6'h1d == cacheLine & 3'h5 == io_addrs[4:2] ? cache_29_line_5 : _GEN_364; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_366 = 6'h1d == cacheLine & 3'h6 == io_addrs[4:2] ? cache_29_line_6 : _GEN_365; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_367 = 6'h1d == cacheLine & 3'h7 == io_addrs[4:2] ? cache_29_line_7 : _GEN_366; // @[Cache.scala 40:{18,18}]
  wire  _GEN_4450 = 6'h1e == cacheLine; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_368 = 6'h1e == cacheLine & 3'h0 == io_addrs[4:2] ? cache_30_line_0 : _GEN_367; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_369 = 6'h1e == cacheLine & 3'h1 == io_addrs[4:2] ? cache_30_line_1 : _GEN_368; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_370 = 6'h1e == cacheLine & 3'h2 == io_addrs[4:2] ? cache_30_line_2 : _GEN_369; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_371 = 6'h1e == cacheLine & 3'h3 == io_addrs[4:2] ? cache_30_line_3 : _GEN_370; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_372 = 6'h1e == cacheLine & 3'h4 == io_addrs[4:2] ? cache_30_line_4 : _GEN_371; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_373 = 6'h1e == cacheLine & 3'h5 == io_addrs[4:2] ? cache_30_line_5 : _GEN_372; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_374 = 6'h1e == cacheLine & 3'h6 == io_addrs[4:2] ? cache_30_line_6 : _GEN_373; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_375 = 6'h1e == cacheLine & 3'h7 == io_addrs[4:2] ? cache_30_line_7 : _GEN_374; // @[Cache.scala 40:{18,18}]
  wire  _GEN_4466 = 6'h1f == cacheLine; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_376 = 6'h1f == cacheLine & 3'h0 == io_addrs[4:2] ? cache_31_line_0 : _GEN_375; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_377 = 6'h1f == cacheLine & 3'h1 == io_addrs[4:2] ? cache_31_line_1 : _GEN_376; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_378 = 6'h1f == cacheLine & 3'h2 == io_addrs[4:2] ? cache_31_line_2 : _GEN_377; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_379 = 6'h1f == cacheLine & 3'h3 == io_addrs[4:2] ? cache_31_line_3 : _GEN_378; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_380 = 6'h1f == cacheLine & 3'h4 == io_addrs[4:2] ? cache_31_line_4 : _GEN_379; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_381 = 6'h1f == cacheLine & 3'h5 == io_addrs[4:2] ? cache_31_line_5 : _GEN_380; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_382 = 6'h1f == cacheLine & 3'h6 == io_addrs[4:2] ? cache_31_line_6 : _GEN_381; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_383 = 6'h1f == cacheLine & 3'h7 == io_addrs[4:2] ? cache_31_line_7 : _GEN_382; // @[Cache.scala 40:{18,18}]
  wire  _GEN_4482 = 6'h20 == cacheLine; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_384 = 6'h20 == cacheLine & 3'h0 == io_addrs[4:2] ? cache_32_line_0 : _GEN_383; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_385 = 6'h20 == cacheLine & 3'h1 == io_addrs[4:2] ? cache_32_line_1 : _GEN_384; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_386 = 6'h20 == cacheLine & 3'h2 == io_addrs[4:2] ? cache_32_line_2 : _GEN_385; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_387 = 6'h20 == cacheLine & 3'h3 == io_addrs[4:2] ? cache_32_line_3 : _GEN_386; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_388 = 6'h20 == cacheLine & 3'h4 == io_addrs[4:2] ? cache_32_line_4 : _GEN_387; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_389 = 6'h20 == cacheLine & 3'h5 == io_addrs[4:2] ? cache_32_line_5 : _GEN_388; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_390 = 6'h20 == cacheLine & 3'h6 == io_addrs[4:2] ? cache_32_line_6 : _GEN_389; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_391 = 6'h20 == cacheLine & 3'h7 == io_addrs[4:2] ? cache_32_line_7 : _GEN_390; // @[Cache.scala 40:{18,18}]
  wire  _GEN_4498 = 6'h21 == cacheLine; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_392 = 6'h21 == cacheLine & 3'h0 == io_addrs[4:2] ? cache_33_line_0 : _GEN_391; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_393 = 6'h21 == cacheLine & 3'h1 == io_addrs[4:2] ? cache_33_line_1 : _GEN_392; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_394 = 6'h21 == cacheLine & 3'h2 == io_addrs[4:2] ? cache_33_line_2 : _GEN_393; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_395 = 6'h21 == cacheLine & 3'h3 == io_addrs[4:2] ? cache_33_line_3 : _GEN_394; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_396 = 6'h21 == cacheLine & 3'h4 == io_addrs[4:2] ? cache_33_line_4 : _GEN_395; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_397 = 6'h21 == cacheLine & 3'h5 == io_addrs[4:2] ? cache_33_line_5 : _GEN_396; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_398 = 6'h21 == cacheLine & 3'h6 == io_addrs[4:2] ? cache_33_line_6 : _GEN_397; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_399 = 6'h21 == cacheLine & 3'h7 == io_addrs[4:2] ? cache_33_line_7 : _GEN_398; // @[Cache.scala 40:{18,18}]
  wire  _GEN_4514 = 6'h22 == cacheLine; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_400 = 6'h22 == cacheLine & 3'h0 == io_addrs[4:2] ? cache_34_line_0 : _GEN_399; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_401 = 6'h22 == cacheLine & 3'h1 == io_addrs[4:2] ? cache_34_line_1 : _GEN_400; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_402 = 6'h22 == cacheLine & 3'h2 == io_addrs[4:2] ? cache_34_line_2 : _GEN_401; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_403 = 6'h22 == cacheLine & 3'h3 == io_addrs[4:2] ? cache_34_line_3 : _GEN_402; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_404 = 6'h22 == cacheLine & 3'h4 == io_addrs[4:2] ? cache_34_line_4 : _GEN_403; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_405 = 6'h22 == cacheLine & 3'h5 == io_addrs[4:2] ? cache_34_line_5 : _GEN_404; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_406 = 6'h22 == cacheLine & 3'h6 == io_addrs[4:2] ? cache_34_line_6 : _GEN_405; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_407 = 6'h22 == cacheLine & 3'h7 == io_addrs[4:2] ? cache_34_line_7 : _GEN_406; // @[Cache.scala 40:{18,18}]
  wire  _GEN_4530 = 6'h23 == cacheLine; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_408 = 6'h23 == cacheLine & 3'h0 == io_addrs[4:2] ? cache_35_line_0 : _GEN_407; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_409 = 6'h23 == cacheLine & 3'h1 == io_addrs[4:2] ? cache_35_line_1 : _GEN_408; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_410 = 6'h23 == cacheLine & 3'h2 == io_addrs[4:2] ? cache_35_line_2 : _GEN_409; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_411 = 6'h23 == cacheLine & 3'h3 == io_addrs[4:2] ? cache_35_line_3 : _GEN_410; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_412 = 6'h23 == cacheLine & 3'h4 == io_addrs[4:2] ? cache_35_line_4 : _GEN_411; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_413 = 6'h23 == cacheLine & 3'h5 == io_addrs[4:2] ? cache_35_line_5 : _GEN_412; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_414 = 6'h23 == cacheLine & 3'h6 == io_addrs[4:2] ? cache_35_line_6 : _GEN_413; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_415 = 6'h23 == cacheLine & 3'h7 == io_addrs[4:2] ? cache_35_line_7 : _GEN_414; // @[Cache.scala 40:{18,18}]
  wire  _GEN_4546 = 6'h24 == cacheLine; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_416 = 6'h24 == cacheLine & 3'h0 == io_addrs[4:2] ? cache_36_line_0 : _GEN_415; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_417 = 6'h24 == cacheLine & 3'h1 == io_addrs[4:2] ? cache_36_line_1 : _GEN_416; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_418 = 6'h24 == cacheLine & 3'h2 == io_addrs[4:2] ? cache_36_line_2 : _GEN_417; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_419 = 6'h24 == cacheLine & 3'h3 == io_addrs[4:2] ? cache_36_line_3 : _GEN_418; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_420 = 6'h24 == cacheLine & 3'h4 == io_addrs[4:2] ? cache_36_line_4 : _GEN_419; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_421 = 6'h24 == cacheLine & 3'h5 == io_addrs[4:2] ? cache_36_line_5 : _GEN_420; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_422 = 6'h24 == cacheLine & 3'h6 == io_addrs[4:2] ? cache_36_line_6 : _GEN_421; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_423 = 6'h24 == cacheLine & 3'h7 == io_addrs[4:2] ? cache_36_line_7 : _GEN_422; // @[Cache.scala 40:{18,18}]
  wire  _GEN_4562 = 6'h25 == cacheLine; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_424 = 6'h25 == cacheLine & 3'h0 == io_addrs[4:2] ? cache_37_line_0 : _GEN_423; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_425 = 6'h25 == cacheLine & 3'h1 == io_addrs[4:2] ? cache_37_line_1 : _GEN_424; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_426 = 6'h25 == cacheLine & 3'h2 == io_addrs[4:2] ? cache_37_line_2 : _GEN_425; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_427 = 6'h25 == cacheLine & 3'h3 == io_addrs[4:2] ? cache_37_line_3 : _GEN_426; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_428 = 6'h25 == cacheLine & 3'h4 == io_addrs[4:2] ? cache_37_line_4 : _GEN_427; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_429 = 6'h25 == cacheLine & 3'h5 == io_addrs[4:2] ? cache_37_line_5 : _GEN_428; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_430 = 6'h25 == cacheLine & 3'h6 == io_addrs[4:2] ? cache_37_line_6 : _GEN_429; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_431 = 6'h25 == cacheLine & 3'h7 == io_addrs[4:2] ? cache_37_line_7 : _GEN_430; // @[Cache.scala 40:{18,18}]
  wire  _GEN_4578 = 6'h26 == cacheLine; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_432 = 6'h26 == cacheLine & 3'h0 == io_addrs[4:2] ? cache_38_line_0 : _GEN_431; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_433 = 6'h26 == cacheLine & 3'h1 == io_addrs[4:2] ? cache_38_line_1 : _GEN_432; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_434 = 6'h26 == cacheLine & 3'h2 == io_addrs[4:2] ? cache_38_line_2 : _GEN_433; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_435 = 6'h26 == cacheLine & 3'h3 == io_addrs[4:2] ? cache_38_line_3 : _GEN_434; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_436 = 6'h26 == cacheLine & 3'h4 == io_addrs[4:2] ? cache_38_line_4 : _GEN_435; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_437 = 6'h26 == cacheLine & 3'h5 == io_addrs[4:2] ? cache_38_line_5 : _GEN_436; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_438 = 6'h26 == cacheLine & 3'h6 == io_addrs[4:2] ? cache_38_line_6 : _GEN_437; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_439 = 6'h26 == cacheLine & 3'h7 == io_addrs[4:2] ? cache_38_line_7 : _GEN_438; // @[Cache.scala 40:{18,18}]
  wire  _GEN_4594 = 6'h27 == cacheLine; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_440 = 6'h27 == cacheLine & 3'h0 == io_addrs[4:2] ? cache_39_line_0 : _GEN_439; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_441 = 6'h27 == cacheLine & 3'h1 == io_addrs[4:2] ? cache_39_line_1 : _GEN_440; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_442 = 6'h27 == cacheLine & 3'h2 == io_addrs[4:2] ? cache_39_line_2 : _GEN_441; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_443 = 6'h27 == cacheLine & 3'h3 == io_addrs[4:2] ? cache_39_line_3 : _GEN_442; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_444 = 6'h27 == cacheLine & 3'h4 == io_addrs[4:2] ? cache_39_line_4 : _GEN_443; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_445 = 6'h27 == cacheLine & 3'h5 == io_addrs[4:2] ? cache_39_line_5 : _GEN_444; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_446 = 6'h27 == cacheLine & 3'h6 == io_addrs[4:2] ? cache_39_line_6 : _GEN_445; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_447 = 6'h27 == cacheLine & 3'h7 == io_addrs[4:2] ? cache_39_line_7 : _GEN_446; // @[Cache.scala 40:{18,18}]
  wire  _GEN_4610 = 6'h28 == cacheLine; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_448 = 6'h28 == cacheLine & 3'h0 == io_addrs[4:2] ? cache_40_line_0 : _GEN_447; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_449 = 6'h28 == cacheLine & 3'h1 == io_addrs[4:2] ? cache_40_line_1 : _GEN_448; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_450 = 6'h28 == cacheLine & 3'h2 == io_addrs[4:2] ? cache_40_line_2 : _GEN_449; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_451 = 6'h28 == cacheLine & 3'h3 == io_addrs[4:2] ? cache_40_line_3 : _GEN_450; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_452 = 6'h28 == cacheLine & 3'h4 == io_addrs[4:2] ? cache_40_line_4 : _GEN_451; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_453 = 6'h28 == cacheLine & 3'h5 == io_addrs[4:2] ? cache_40_line_5 : _GEN_452; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_454 = 6'h28 == cacheLine & 3'h6 == io_addrs[4:2] ? cache_40_line_6 : _GEN_453; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_455 = 6'h28 == cacheLine & 3'h7 == io_addrs[4:2] ? cache_40_line_7 : _GEN_454; // @[Cache.scala 40:{18,18}]
  wire  _GEN_4626 = 6'h29 == cacheLine; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_456 = 6'h29 == cacheLine & 3'h0 == io_addrs[4:2] ? cache_41_line_0 : _GEN_455; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_457 = 6'h29 == cacheLine & 3'h1 == io_addrs[4:2] ? cache_41_line_1 : _GEN_456; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_458 = 6'h29 == cacheLine & 3'h2 == io_addrs[4:2] ? cache_41_line_2 : _GEN_457; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_459 = 6'h29 == cacheLine & 3'h3 == io_addrs[4:2] ? cache_41_line_3 : _GEN_458; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_460 = 6'h29 == cacheLine & 3'h4 == io_addrs[4:2] ? cache_41_line_4 : _GEN_459; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_461 = 6'h29 == cacheLine & 3'h5 == io_addrs[4:2] ? cache_41_line_5 : _GEN_460; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_462 = 6'h29 == cacheLine & 3'h6 == io_addrs[4:2] ? cache_41_line_6 : _GEN_461; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_463 = 6'h29 == cacheLine & 3'h7 == io_addrs[4:2] ? cache_41_line_7 : _GEN_462; // @[Cache.scala 40:{18,18}]
  wire  _GEN_4642 = 6'h2a == cacheLine; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_464 = 6'h2a == cacheLine & 3'h0 == io_addrs[4:2] ? cache_42_line_0 : _GEN_463; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_465 = 6'h2a == cacheLine & 3'h1 == io_addrs[4:2] ? cache_42_line_1 : _GEN_464; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_466 = 6'h2a == cacheLine & 3'h2 == io_addrs[4:2] ? cache_42_line_2 : _GEN_465; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_467 = 6'h2a == cacheLine & 3'h3 == io_addrs[4:2] ? cache_42_line_3 : _GEN_466; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_468 = 6'h2a == cacheLine & 3'h4 == io_addrs[4:2] ? cache_42_line_4 : _GEN_467; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_469 = 6'h2a == cacheLine & 3'h5 == io_addrs[4:2] ? cache_42_line_5 : _GEN_468; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_470 = 6'h2a == cacheLine & 3'h6 == io_addrs[4:2] ? cache_42_line_6 : _GEN_469; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_471 = 6'h2a == cacheLine & 3'h7 == io_addrs[4:2] ? cache_42_line_7 : _GEN_470; // @[Cache.scala 40:{18,18}]
  wire  _GEN_4658 = 6'h2b == cacheLine; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_472 = 6'h2b == cacheLine & 3'h0 == io_addrs[4:2] ? cache_43_line_0 : _GEN_471; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_473 = 6'h2b == cacheLine & 3'h1 == io_addrs[4:2] ? cache_43_line_1 : _GEN_472; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_474 = 6'h2b == cacheLine & 3'h2 == io_addrs[4:2] ? cache_43_line_2 : _GEN_473; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_475 = 6'h2b == cacheLine & 3'h3 == io_addrs[4:2] ? cache_43_line_3 : _GEN_474; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_476 = 6'h2b == cacheLine & 3'h4 == io_addrs[4:2] ? cache_43_line_4 : _GEN_475; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_477 = 6'h2b == cacheLine & 3'h5 == io_addrs[4:2] ? cache_43_line_5 : _GEN_476; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_478 = 6'h2b == cacheLine & 3'h6 == io_addrs[4:2] ? cache_43_line_6 : _GEN_477; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_479 = 6'h2b == cacheLine & 3'h7 == io_addrs[4:2] ? cache_43_line_7 : _GEN_478; // @[Cache.scala 40:{18,18}]
  wire  _GEN_4674 = 6'h2c == cacheLine; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_480 = 6'h2c == cacheLine & 3'h0 == io_addrs[4:2] ? cache_44_line_0 : _GEN_479; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_481 = 6'h2c == cacheLine & 3'h1 == io_addrs[4:2] ? cache_44_line_1 : _GEN_480; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_482 = 6'h2c == cacheLine & 3'h2 == io_addrs[4:2] ? cache_44_line_2 : _GEN_481; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_483 = 6'h2c == cacheLine & 3'h3 == io_addrs[4:2] ? cache_44_line_3 : _GEN_482; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_484 = 6'h2c == cacheLine & 3'h4 == io_addrs[4:2] ? cache_44_line_4 : _GEN_483; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_485 = 6'h2c == cacheLine & 3'h5 == io_addrs[4:2] ? cache_44_line_5 : _GEN_484; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_486 = 6'h2c == cacheLine & 3'h6 == io_addrs[4:2] ? cache_44_line_6 : _GEN_485; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_487 = 6'h2c == cacheLine & 3'h7 == io_addrs[4:2] ? cache_44_line_7 : _GEN_486; // @[Cache.scala 40:{18,18}]
  wire  _GEN_4690 = 6'h2d == cacheLine; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_488 = 6'h2d == cacheLine & 3'h0 == io_addrs[4:2] ? cache_45_line_0 : _GEN_487; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_489 = 6'h2d == cacheLine & 3'h1 == io_addrs[4:2] ? cache_45_line_1 : _GEN_488; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_490 = 6'h2d == cacheLine & 3'h2 == io_addrs[4:2] ? cache_45_line_2 : _GEN_489; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_491 = 6'h2d == cacheLine & 3'h3 == io_addrs[4:2] ? cache_45_line_3 : _GEN_490; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_492 = 6'h2d == cacheLine & 3'h4 == io_addrs[4:2] ? cache_45_line_4 : _GEN_491; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_493 = 6'h2d == cacheLine & 3'h5 == io_addrs[4:2] ? cache_45_line_5 : _GEN_492; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_494 = 6'h2d == cacheLine & 3'h6 == io_addrs[4:2] ? cache_45_line_6 : _GEN_493; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_495 = 6'h2d == cacheLine & 3'h7 == io_addrs[4:2] ? cache_45_line_7 : _GEN_494; // @[Cache.scala 40:{18,18}]
  wire  _GEN_4706 = 6'h2e == cacheLine; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_496 = 6'h2e == cacheLine & 3'h0 == io_addrs[4:2] ? cache_46_line_0 : _GEN_495; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_497 = 6'h2e == cacheLine & 3'h1 == io_addrs[4:2] ? cache_46_line_1 : _GEN_496; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_498 = 6'h2e == cacheLine & 3'h2 == io_addrs[4:2] ? cache_46_line_2 : _GEN_497; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_499 = 6'h2e == cacheLine & 3'h3 == io_addrs[4:2] ? cache_46_line_3 : _GEN_498; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_500 = 6'h2e == cacheLine & 3'h4 == io_addrs[4:2] ? cache_46_line_4 : _GEN_499; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_501 = 6'h2e == cacheLine & 3'h5 == io_addrs[4:2] ? cache_46_line_5 : _GEN_500; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_502 = 6'h2e == cacheLine & 3'h6 == io_addrs[4:2] ? cache_46_line_6 : _GEN_501; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_503 = 6'h2e == cacheLine & 3'h7 == io_addrs[4:2] ? cache_46_line_7 : _GEN_502; // @[Cache.scala 40:{18,18}]
  wire  _GEN_4722 = 6'h2f == cacheLine; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_504 = 6'h2f == cacheLine & 3'h0 == io_addrs[4:2] ? cache_47_line_0 : _GEN_503; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_505 = 6'h2f == cacheLine & 3'h1 == io_addrs[4:2] ? cache_47_line_1 : _GEN_504; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_506 = 6'h2f == cacheLine & 3'h2 == io_addrs[4:2] ? cache_47_line_2 : _GEN_505; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_507 = 6'h2f == cacheLine & 3'h3 == io_addrs[4:2] ? cache_47_line_3 : _GEN_506; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_508 = 6'h2f == cacheLine & 3'h4 == io_addrs[4:2] ? cache_47_line_4 : _GEN_507; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_509 = 6'h2f == cacheLine & 3'h5 == io_addrs[4:2] ? cache_47_line_5 : _GEN_508; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_510 = 6'h2f == cacheLine & 3'h6 == io_addrs[4:2] ? cache_47_line_6 : _GEN_509; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_511 = 6'h2f == cacheLine & 3'h7 == io_addrs[4:2] ? cache_47_line_7 : _GEN_510; // @[Cache.scala 40:{18,18}]
  wire  _GEN_4738 = 6'h30 == cacheLine; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_512 = 6'h30 == cacheLine & 3'h0 == io_addrs[4:2] ? cache_48_line_0 : _GEN_511; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_513 = 6'h30 == cacheLine & 3'h1 == io_addrs[4:2] ? cache_48_line_1 : _GEN_512; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_514 = 6'h30 == cacheLine & 3'h2 == io_addrs[4:2] ? cache_48_line_2 : _GEN_513; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_515 = 6'h30 == cacheLine & 3'h3 == io_addrs[4:2] ? cache_48_line_3 : _GEN_514; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_516 = 6'h30 == cacheLine & 3'h4 == io_addrs[4:2] ? cache_48_line_4 : _GEN_515; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_517 = 6'h30 == cacheLine & 3'h5 == io_addrs[4:2] ? cache_48_line_5 : _GEN_516; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_518 = 6'h30 == cacheLine & 3'h6 == io_addrs[4:2] ? cache_48_line_6 : _GEN_517; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_519 = 6'h30 == cacheLine & 3'h7 == io_addrs[4:2] ? cache_48_line_7 : _GEN_518; // @[Cache.scala 40:{18,18}]
  wire  _GEN_4754 = 6'h31 == cacheLine; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_520 = 6'h31 == cacheLine & 3'h0 == io_addrs[4:2] ? cache_49_line_0 : _GEN_519; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_521 = 6'h31 == cacheLine & 3'h1 == io_addrs[4:2] ? cache_49_line_1 : _GEN_520; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_522 = 6'h31 == cacheLine & 3'h2 == io_addrs[4:2] ? cache_49_line_2 : _GEN_521; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_523 = 6'h31 == cacheLine & 3'h3 == io_addrs[4:2] ? cache_49_line_3 : _GEN_522; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_524 = 6'h31 == cacheLine & 3'h4 == io_addrs[4:2] ? cache_49_line_4 : _GEN_523; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_525 = 6'h31 == cacheLine & 3'h5 == io_addrs[4:2] ? cache_49_line_5 : _GEN_524; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_526 = 6'h31 == cacheLine & 3'h6 == io_addrs[4:2] ? cache_49_line_6 : _GEN_525; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_527 = 6'h31 == cacheLine & 3'h7 == io_addrs[4:2] ? cache_49_line_7 : _GEN_526; // @[Cache.scala 40:{18,18}]
  wire  _GEN_4770 = 6'h32 == cacheLine; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_528 = 6'h32 == cacheLine & 3'h0 == io_addrs[4:2] ? cache_50_line_0 : _GEN_527; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_529 = 6'h32 == cacheLine & 3'h1 == io_addrs[4:2] ? cache_50_line_1 : _GEN_528; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_530 = 6'h32 == cacheLine & 3'h2 == io_addrs[4:2] ? cache_50_line_2 : _GEN_529; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_531 = 6'h32 == cacheLine & 3'h3 == io_addrs[4:2] ? cache_50_line_3 : _GEN_530; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_532 = 6'h32 == cacheLine & 3'h4 == io_addrs[4:2] ? cache_50_line_4 : _GEN_531; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_533 = 6'h32 == cacheLine & 3'h5 == io_addrs[4:2] ? cache_50_line_5 : _GEN_532; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_534 = 6'h32 == cacheLine & 3'h6 == io_addrs[4:2] ? cache_50_line_6 : _GEN_533; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_535 = 6'h32 == cacheLine & 3'h7 == io_addrs[4:2] ? cache_50_line_7 : _GEN_534; // @[Cache.scala 40:{18,18}]
  wire  _GEN_4786 = 6'h33 == cacheLine; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_536 = 6'h33 == cacheLine & 3'h0 == io_addrs[4:2] ? cache_51_line_0 : _GEN_535; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_537 = 6'h33 == cacheLine & 3'h1 == io_addrs[4:2] ? cache_51_line_1 : _GEN_536; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_538 = 6'h33 == cacheLine & 3'h2 == io_addrs[4:2] ? cache_51_line_2 : _GEN_537; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_539 = 6'h33 == cacheLine & 3'h3 == io_addrs[4:2] ? cache_51_line_3 : _GEN_538; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_540 = 6'h33 == cacheLine & 3'h4 == io_addrs[4:2] ? cache_51_line_4 : _GEN_539; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_541 = 6'h33 == cacheLine & 3'h5 == io_addrs[4:2] ? cache_51_line_5 : _GEN_540; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_542 = 6'h33 == cacheLine & 3'h6 == io_addrs[4:2] ? cache_51_line_6 : _GEN_541; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_543 = 6'h33 == cacheLine & 3'h7 == io_addrs[4:2] ? cache_51_line_7 : _GEN_542; // @[Cache.scala 40:{18,18}]
  wire  _GEN_4802 = 6'h34 == cacheLine; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_544 = 6'h34 == cacheLine & 3'h0 == io_addrs[4:2] ? cache_52_line_0 : _GEN_543; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_545 = 6'h34 == cacheLine & 3'h1 == io_addrs[4:2] ? cache_52_line_1 : _GEN_544; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_546 = 6'h34 == cacheLine & 3'h2 == io_addrs[4:2] ? cache_52_line_2 : _GEN_545; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_547 = 6'h34 == cacheLine & 3'h3 == io_addrs[4:2] ? cache_52_line_3 : _GEN_546; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_548 = 6'h34 == cacheLine & 3'h4 == io_addrs[4:2] ? cache_52_line_4 : _GEN_547; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_549 = 6'h34 == cacheLine & 3'h5 == io_addrs[4:2] ? cache_52_line_5 : _GEN_548; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_550 = 6'h34 == cacheLine & 3'h6 == io_addrs[4:2] ? cache_52_line_6 : _GEN_549; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_551 = 6'h34 == cacheLine & 3'h7 == io_addrs[4:2] ? cache_52_line_7 : _GEN_550; // @[Cache.scala 40:{18,18}]
  wire  _GEN_4818 = 6'h35 == cacheLine; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_552 = 6'h35 == cacheLine & 3'h0 == io_addrs[4:2] ? cache_53_line_0 : _GEN_551; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_553 = 6'h35 == cacheLine & 3'h1 == io_addrs[4:2] ? cache_53_line_1 : _GEN_552; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_554 = 6'h35 == cacheLine & 3'h2 == io_addrs[4:2] ? cache_53_line_2 : _GEN_553; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_555 = 6'h35 == cacheLine & 3'h3 == io_addrs[4:2] ? cache_53_line_3 : _GEN_554; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_556 = 6'h35 == cacheLine & 3'h4 == io_addrs[4:2] ? cache_53_line_4 : _GEN_555; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_557 = 6'h35 == cacheLine & 3'h5 == io_addrs[4:2] ? cache_53_line_5 : _GEN_556; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_558 = 6'h35 == cacheLine & 3'h6 == io_addrs[4:2] ? cache_53_line_6 : _GEN_557; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_559 = 6'h35 == cacheLine & 3'h7 == io_addrs[4:2] ? cache_53_line_7 : _GEN_558; // @[Cache.scala 40:{18,18}]
  wire  _GEN_4834 = 6'h36 == cacheLine; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_560 = 6'h36 == cacheLine & 3'h0 == io_addrs[4:2] ? cache_54_line_0 : _GEN_559; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_561 = 6'h36 == cacheLine & 3'h1 == io_addrs[4:2] ? cache_54_line_1 : _GEN_560; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_562 = 6'h36 == cacheLine & 3'h2 == io_addrs[4:2] ? cache_54_line_2 : _GEN_561; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_563 = 6'h36 == cacheLine & 3'h3 == io_addrs[4:2] ? cache_54_line_3 : _GEN_562; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_564 = 6'h36 == cacheLine & 3'h4 == io_addrs[4:2] ? cache_54_line_4 : _GEN_563; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_565 = 6'h36 == cacheLine & 3'h5 == io_addrs[4:2] ? cache_54_line_5 : _GEN_564; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_566 = 6'h36 == cacheLine & 3'h6 == io_addrs[4:2] ? cache_54_line_6 : _GEN_565; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_567 = 6'h36 == cacheLine & 3'h7 == io_addrs[4:2] ? cache_54_line_7 : _GEN_566; // @[Cache.scala 40:{18,18}]
  wire  _GEN_4850 = 6'h37 == cacheLine; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_568 = 6'h37 == cacheLine & 3'h0 == io_addrs[4:2] ? cache_55_line_0 : _GEN_567; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_569 = 6'h37 == cacheLine & 3'h1 == io_addrs[4:2] ? cache_55_line_1 : _GEN_568; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_570 = 6'h37 == cacheLine & 3'h2 == io_addrs[4:2] ? cache_55_line_2 : _GEN_569; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_571 = 6'h37 == cacheLine & 3'h3 == io_addrs[4:2] ? cache_55_line_3 : _GEN_570; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_572 = 6'h37 == cacheLine & 3'h4 == io_addrs[4:2] ? cache_55_line_4 : _GEN_571; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_573 = 6'h37 == cacheLine & 3'h5 == io_addrs[4:2] ? cache_55_line_5 : _GEN_572; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_574 = 6'h37 == cacheLine & 3'h6 == io_addrs[4:2] ? cache_55_line_6 : _GEN_573; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_575 = 6'h37 == cacheLine & 3'h7 == io_addrs[4:2] ? cache_55_line_7 : _GEN_574; // @[Cache.scala 40:{18,18}]
  wire  _GEN_4866 = 6'h38 == cacheLine; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_576 = 6'h38 == cacheLine & 3'h0 == io_addrs[4:2] ? cache_56_line_0 : _GEN_575; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_577 = 6'h38 == cacheLine & 3'h1 == io_addrs[4:2] ? cache_56_line_1 : _GEN_576; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_578 = 6'h38 == cacheLine & 3'h2 == io_addrs[4:2] ? cache_56_line_2 : _GEN_577; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_579 = 6'h38 == cacheLine & 3'h3 == io_addrs[4:2] ? cache_56_line_3 : _GEN_578; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_580 = 6'h38 == cacheLine & 3'h4 == io_addrs[4:2] ? cache_56_line_4 : _GEN_579; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_581 = 6'h38 == cacheLine & 3'h5 == io_addrs[4:2] ? cache_56_line_5 : _GEN_580; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_582 = 6'h38 == cacheLine & 3'h6 == io_addrs[4:2] ? cache_56_line_6 : _GEN_581; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_583 = 6'h38 == cacheLine & 3'h7 == io_addrs[4:2] ? cache_56_line_7 : _GEN_582; // @[Cache.scala 40:{18,18}]
  wire  _GEN_4882 = 6'h39 == cacheLine; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_584 = 6'h39 == cacheLine & 3'h0 == io_addrs[4:2] ? cache_57_line_0 : _GEN_583; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_585 = 6'h39 == cacheLine & 3'h1 == io_addrs[4:2] ? cache_57_line_1 : _GEN_584; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_586 = 6'h39 == cacheLine & 3'h2 == io_addrs[4:2] ? cache_57_line_2 : _GEN_585; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_587 = 6'h39 == cacheLine & 3'h3 == io_addrs[4:2] ? cache_57_line_3 : _GEN_586; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_588 = 6'h39 == cacheLine & 3'h4 == io_addrs[4:2] ? cache_57_line_4 : _GEN_587; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_589 = 6'h39 == cacheLine & 3'h5 == io_addrs[4:2] ? cache_57_line_5 : _GEN_588; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_590 = 6'h39 == cacheLine & 3'h6 == io_addrs[4:2] ? cache_57_line_6 : _GEN_589; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_591 = 6'h39 == cacheLine & 3'h7 == io_addrs[4:2] ? cache_57_line_7 : _GEN_590; // @[Cache.scala 40:{18,18}]
  wire  _GEN_4898 = 6'h3a == cacheLine; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_592 = 6'h3a == cacheLine & 3'h0 == io_addrs[4:2] ? cache_58_line_0 : _GEN_591; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_593 = 6'h3a == cacheLine & 3'h1 == io_addrs[4:2] ? cache_58_line_1 : _GEN_592; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_594 = 6'h3a == cacheLine & 3'h2 == io_addrs[4:2] ? cache_58_line_2 : _GEN_593; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_595 = 6'h3a == cacheLine & 3'h3 == io_addrs[4:2] ? cache_58_line_3 : _GEN_594; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_596 = 6'h3a == cacheLine & 3'h4 == io_addrs[4:2] ? cache_58_line_4 : _GEN_595; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_597 = 6'h3a == cacheLine & 3'h5 == io_addrs[4:2] ? cache_58_line_5 : _GEN_596; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_598 = 6'h3a == cacheLine & 3'h6 == io_addrs[4:2] ? cache_58_line_6 : _GEN_597; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_599 = 6'h3a == cacheLine & 3'h7 == io_addrs[4:2] ? cache_58_line_7 : _GEN_598; // @[Cache.scala 40:{18,18}]
  wire  _GEN_4914 = 6'h3b == cacheLine; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_600 = 6'h3b == cacheLine & 3'h0 == io_addrs[4:2] ? cache_59_line_0 : _GEN_599; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_601 = 6'h3b == cacheLine & 3'h1 == io_addrs[4:2] ? cache_59_line_1 : _GEN_600; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_602 = 6'h3b == cacheLine & 3'h2 == io_addrs[4:2] ? cache_59_line_2 : _GEN_601; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_603 = 6'h3b == cacheLine & 3'h3 == io_addrs[4:2] ? cache_59_line_3 : _GEN_602; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_604 = 6'h3b == cacheLine & 3'h4 == io_addrs[4:2] ? cache_59_line_4 : _GEN_603; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_605 = 6'h3b == cacheLine & 3'h5 == io_addrs[4:2] ? cache_59_line_5 : _GEN_604; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_606 = 6'h3b == cacheLine & 3'h6 == io_addrs[4:2] ? cache_59_line_6 : _GEN_605; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_607 = 6'h3b == cacheLine & 3'h7 == io_addrs[4:2] ? cache_59_line_7 : _GEN_606; // @[Cache.scala 40:{18,18}]
  wire  _GEN_4930 = 6'h3c == cacheLine; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_608 = 6'h3c == cacheLine & 3'h0 == io_addrs[4:2] ? cache_60_line_0 : _GEN_607; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_609 = 6'h3c == cacheLine & 3'h1 == io_addrs[4:2] ? cache_60_line_1 : _GEN_608; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_610 = 6'h3c == cacheLine & 3'h2 == io_addrs[4:2] ? cache_60_line_2 : _GEN_609; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_611 = 6'h3c == cacheLine & 3'h3 == io_addrs[4:2] ? cache_60_line_3 : _GEN_610; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_612 = 6'h3c == cacheLine & 3'h4 == io_addrs[4:2] ? cache_60_line_4 : _GEN_611; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_613 = 6'h3c == cacheLine & 3'h5 == io_addrs[4:2] ? cache_60_line_5 : _GEN_612; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_614 = 6'h3c == cacheLine & 3'h6 == io_addrs[4:2] ? cache_60_line_6 : _GEN_613; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_615 = 6'h3c == cacheLine & 3'h7 == io_addrs[4:2] ? cache_60_line_7 : _GEN_614; // @[Cache.scala 40:{18,18}]
  wire  _GEN_4946 = 6'h3d == cacheLine; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_616 = 6'h3d == cacheLine & 3'h0 == io_addrs[4:2] ? cache_61_line_0 : _GEN_615; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_617 = 6'h3d == cacheLine & 3'h1 == io_addrs[4:2] ? cache_61_line_1 : _GEN_616; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_618 = 6'h3d == cacheLine & 3'h2 == io_addrs[4:2] ? cache_61_line_2 : _GEN_617; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_619 = 6'h3d == cacheLine & 3'h3 == io_addrs[4:2] ? cache_61_line_3 : _GEN_618; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_620 = 6'h3d == cacheLine & 3'h4 == io_addrs[4:2] ? cache_61_line_4 : _GEN_619; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_621 = 6'h3d == cacheLine & 3'h5 == io_addrs[4:2] ? cache_61_line_5 : _GEN_620; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_622 = 6'h3d == cacheLine & 3'h6 == io_addrs[4:2] ? cache_61_line_6 : _GEN_621; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_623 = 6'h3d == cacheLine & 3'h7 == io_addrs[4:2] ? cache_61_line_7 : _GEN_622; // @[Cache.scala 40:{18,18}]
  wire  _GEN_4962 = 6'h3e == cacheLine; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_624 = 6'h3e == cacheLine & 3'h0 == io_addrs[4:2] ? cache_62_line_0 : _GEN_623; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_625 = 6'h3e == cacheLine & 3'h1 == io_addrs[4:2] ? cache_62_line_1 : _GEN_624; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_626 = 6'h3e == cacheLine & 3'h2 == io_addrs[4:2] ? cache_62_line_2 : _GEN_625; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_627 = 6'h3e == cacheLine & 3'h3 == io_addrs[4:2] ? cache_62_line_3 : _GEN_626; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_628 = 6'h3e == cacheLine & 3'h4 == io_addrs[4:2] ? cache_62_line_4 : _GEN_627; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_629 = 6'h3e == cacheLine & 3'h5 == io_addrs[4:2] ? cache_62_line_5 : _GEN_628; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_630 = 6'h3e == cacheLine & 3'h6 == io_addrs[4:2] ? cache_62_line_6 : _GEN_629; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_631 = 6'h3e == cacheLine & 3'h7 == io_addrs[4:2] ? cache_62_line_7 : _GEN_630; // @[Cache.scala 40:{18,18}]
  wire  _GEN_4978 = 6'h3f == cacheLine; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_632 = 6'h3f == cacheLine & 3'h0 == io_addrs[4:2] ? cache_63_line_0 : _GEN_631; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_633 = 6'h3f == cacheLine & 3'h1 == io_addrs[4:2] ? cache_63_line_1 : _GEN_632; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_634 = 6'h3f == cacheLine & 3'h2 == io_addrs[4:2] ? cache_63_line_2 : _GEN_633; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_635 = 6'h3f == cacheLine & 3'h3 == io_addrs[4:2] ? cache_63_line_3 : _GEN_634; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_636 = 6'h3f == cacheLine & 3'h4 == io_addrs[4:2] ? cache_63_line_4 : _GEN_635; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_637 = 6'h3f == cacheLine & 3'h5 == io_addrs[4:2] ? cache_63_line_5 : _GEN_636; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_638 = 6'h3f == cacheLine & 3'h6 == io_addrs[4:2] ? cache_63_line_6 : _GEN_637; // @[Cache.scala 40:{18,18}]
  wire [31:0] _GEN_639 = 6'h3f == cacheLine & 3'h7 == io_addrs[4:2] ? cache_63_line_7 : _GEN_638; // @[Cache.scala 40:{18,18}]
  wire [10:0] _addrsBuffer_T = {_GEN_127,cacheLine}; // @[Cache.scala 44:39]
  wire [31:0] _GEN_641 = 6'h1 == cacheLine ? cache_1_line_1 : cache_0_line_1; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_642 = 6'h2 == cacheLine ? cache_2_line_1 : _GEN_641; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_643 = 6'h3 == cacheLine ? cache_3_line_1 : _GEN_642; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_644 = 6'h4 == cacheLine ? cache_4_line_1 : _GEN_643; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_645 = 6'h5 == cacheLine ? cache_5_line_1 : _GEN_644; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_646 = 6'h6 == cacheLine ? cache_6_line_1 : _GEN_645; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_647 = 6'h7 == cacheLine ? cache_7_line_1 : _GEN_646; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_648 = 6'h8 == cacheLine ? cache_8_line_1 : _GEN_647; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_649 = 6'h9 == cacheLine ? cache_9_line_1 : _GEN_648; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_650 = 6'ha == cacheLine ? cache_10_line_1 : _GEN_649; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_651 = 6'hb == cacheLine ? cache_11_line_1 : _GEN_650; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_652 = 6'hc == cacheLine ? cache_12_line_1 : _GEN_651; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_653 = 6'hd == cacheLine ? cache_13_line_1 : _GEN_652; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_654 = 6'he == cacheLine ? cache_14_line_1 : _GEN_653; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_655 = 6'hf == cacheLine ? cache_15_line_1 : _GEN_654; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_656 = 6'h10 == cacheLine ? cache_16_line_1 : _GEN_655; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_657 = 6'h11 == cacheLine ? cache_17_line_1 : _GEN_656; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_658 = 6'h12 == cacheLine ? cache_18_line_1 : _GEN_657; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_659 = 6'h13 == cacheLine ? cache_19_line_1 : _GEN_658; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_660 = 6'h14 == cacheLine ? cache_20_line_1 : _GEN_659; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_661 = 6'h15 == cacheLine ? cache_21_line_1 : _GEN_660; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_662 = 6'h16 == cacheLine ? cache_22_line_1 : _GEN_661; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_663 = 6'h17 == cacheLine ? cache_23_line_1 : _GEN_662; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_664 = 6'h18 == cacheLine ? cache_24_line_1 : _GEN_663; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_665 = 6'h19 == cacheLine ? cache_25_line_1 : _GEN_664; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_666 = 6'h1a == cacheLine ? cache_26_line_1 : _GEN_665; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_667 = 6'h1b == cacheLine ? cache_27_line_1 : _GEN_666; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_668 = 6'h1c == cacheLine ? cache_28_line_1 : _GEN_667; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_669 = 6'h1d == cacheLine ? cache_29_line_1 : _GEN_668; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_670 = 6'h1e == cacheLine ? cache_30_line_1 : _GEN_669; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_671 = 6'h1f == cacheLine ? cache_31_line_1 : _GEN_670; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_672 = 6'h20 == cacheLine ? cache_32_line_1 : _GEN_671; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_673 = 6'h21 == cacheLine ? cache_33_line_1 : _GEN_672; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_674 = 6'h22 == cacheLine ? cache_34_line_1 : _GEN_673; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_675 = 6'h23 == cacheLine ? cache_35_line_1 : _GEN_674; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_676 = 6'h24 == cacheLine ? cache_36_line_1 : _GEN_675; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_677 = 6'h25 == cacheLine ? cache_37_line_1 : _GEN_676; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_678 = 6'h26 == cacheLine ? cache_38_line_1 : _GEN_677; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_679 = 6'h27 == cacheLine ? cache_39_line_1 : _GEN_678; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_680 = 6'h28 == cacheLine ? cache_40_line_1 : _GEN_679; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_681 = 6'h29 == cacheLine ? cache_41_line_1 : _GEN_680; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_682 = 6'h2a == cacheLine ? cache_42_line_1 : _GEN_681; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_683 = 6'h2b == cacheLine ? cache_43_line_1 : _GEN_682; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_684 = 6'h2c == cacheLine ? cache_44_line_1 : _GEN_683; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_685 = 6'h2d == cacheLine ? cache_45_line_1 : _GEN_684; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_686 = 6'h2e == cacheLine ? cache_46_line_1 : _GEN_685; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_687 = 6'h2f == cacheLine ? cache_47_line_1 : _GEN_686; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_688 = 6'h30 == cacheLine ? cache_48_line_1 : _GEN_687; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_689 = 6'h31 == cacheLine ? cache_49_line_1 : _GEN_688; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_690 = 6'h32 == cacheLine ? cache_50_line_1 : _GEN_689; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_691 = 6'h33 == cacheLine ? cache_51_line_1 : _GEN_690; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_692 = 6'h34 == cacheLine ? cache_52_line_1 : _GEN_691; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_693 = 6'h35 == cacheLine ? cache_53_line_1 : _GEN_692; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_694 = 6'h36 == cacheLine ? cache_54_line_1 : _GEN_693; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_695 = 6'h37 == cacheLine ? cache_55_line_1 : _GEN_694; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_696 = 6'h38 == cacheLine ? cache_56_line_1 : _GEN_695; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_697 = 6'h39 == cacheLine ? cache_57_line_1 : _GEN_696; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_698 = 6'h3a == cacheLine ? cache_58_line_1 : _GEN_697; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_699 = 6'h3b == cacheLine ? cache_59_line_1 : _GEN_698; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_700 = 6'h3c == cacheLine ? cache_60_line_1 : _GEN_699; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_701 = 6'h3d == cacheLine ? cache_61_line_1 : _GEN_700; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_702 = 6'h3e == cacheLine ? cache_62_line_1 : _GEN_701; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_703 = 6'h3f == cacheLine ? cache_63_line_1 : _GEN_702; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_705 = 6'h1 == cacheLine ? cache_1_line_0 : cache_0_line_0; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_706 = 6'h2 == cacheLine ? cache_2_line_0 : _GEN_705; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_707 = 6'h3 == cacheLine ? cache_3_line_0 : _GEN_706; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_708 = 6'h4 == cacheLine ? cache_4_line_0 : _GEN_707; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_709 = 6'h5 == cacheLine ? cache_5_line_0 : _GEN_708; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_710 = 6'h6 == cacheLine ? cache_6_line_0 : _GEN_709; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_711 = 6'h7 == cacheLine ? cache_7_line_0 : _GEN_710; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_712 = 6'h8 == cacheLine ? cache_8_line_0 : _GEN_711; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_713 = 6'h9 == cacheLine ? cache_9_line_0 : _GEN_712; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_714 = 6'ha == cacheLine ? cache_10_line_0 : _GEN_713; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_715 = 6'hb == cacheLine ? cache_11_line_0 : _GEN_714; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_716 = 6'hc == cacheLine ? cache_12_line_0 : _GEN_715; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_717 = 6'hd == cacheLine ? cache_13_line_0 : _GEN_716; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_718 = 6'he == cacheLine ? cache_14_line_0 : _GEN_717; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_719 = 6'hf == cacheLine ? cache_15_line_0 : _GEN_718; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_720 = 6'h10 == cacheLine ? cache_16_line_0 : _GEN_719; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_721 = 6'h11 == cacheLine ? cache_17_line_0 : _GEN_720; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_722 = 6'h12 == cacheLine ? cache_18_line_0 : _GEN_721; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_723 = 6'h13 == cacheLine ? cache_19_line_0 : _GEN_722; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_724 = 6'h14 == cacheLine ? cache_20_line_0 : _GEN_723; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_725 = 6'h15 == cacheLine ? cache_21_line_0 : _GEN_724; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_726 = 6'h16 == cacheLine ? cache_22_line_0 : _GEN_725; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_727 = 6'h17 == cacheLine ? cache_23_line_0 : _GEN_726; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_728 = 6'h18 == cacheLine ? cache_24_line_0 : _GEN_727; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_729 = 6'h19 == cacheLine ? cache_25_line_0 : _GEN_728; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_730 = 6'h1a == cacheLine ? cache_26_line_0 : _GEN_729; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_731 = 6'h1b == cacheLine ? cache_27_line_0 : _GEN_730; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_732 = 6'h1c == cacheLine ? cache_28_line_0 : _GEN_731; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_733 = 6'h1d == cacheLine ? cache_29_line_0 : _GEN_732; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_734 = 6'h1e == cacheLine ? cache_30_line_0 : _GEN_733; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_735 = 6'h1f == cacheLine ? cache_31_line_0 : _GEN_734; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_736 = 6'h20 == cacheLine ? cache_32_line_0 : _GEN_735; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_737 = 6'h21 == cacheLine ? cache_33_line_0 : _GEN_736; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_738 = 6'h22 == cacheLine ? cache_34_line_0 : _GEN_737; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_739 = 6'h23 == cacheLine ? cache_35_line_0 : _GEN_738; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_740 = 6'h24 == cacheLine ? cache_36_line_0 : _GEN_739; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_741 = 6'h25 == cacheLine ? cache_37_line_0 : _GEN_740; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_742 = 6'h26 == cacheLine ? cache_38_line_0 : _GEN_741; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_743 = 6'h27 == cacheLine ? cache_39_line_0 : _GEN_742; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_744 = 6'h28 == cacheLine ? cache_40_line_0 : _GEN_743; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_745 = 6'h29 == cacheLine ? cache_41_line_0 : _GEN_744; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_746 = 6'h2a == cacheLine ? cache_42_line_0 : _GEN_745; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_747 = 6'h2b == cacheLine ? cache_43_line_0 : _GEN_746; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_748 = 6'h2c == cacheLine ? cache_44_line_0 : _GEN_747; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_749 = 6'h2d == cacheLine ? cache_45_line_0 : _GEN_748; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_750 = 6'h2e == cacheLine ? cache_46_line_0 : _GEN_749; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_751 = 6'h2f == cacheLine ? cache_47_line_0 : _GEN_750; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_752 = 6'h30 == cacheLine ? cache_48_line_0 : _GEN_751; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_753 = 6'h31 == cacheLine ? cache_49_line_0 : _GEN_752; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_754 = 6'h32 == cacheLine ? cache_50_line_0 : _GEN_753; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_755 = 6'h33 == cacheLine ? cache_51_line_0 : _GEN_754; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_756 = 6'h34 == cacheLine ? cache_52_line_0 : _GEN_755; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_757 = 6'h35 == cacheLine ? cache_53_line_0 : _GEN_756; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_758 = 6'h36 == cacheLine ? cache_54_line_0 : _GEN_757; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_759 = 6'h37 == cacheLine ? cache_55_line_0 : _GEN_758; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_760 = 6'h38 == cacheLine ? cache_56_line_0 : _GEN_759; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_761 = 6'h39 == cacheLine ? cache_57_line_0 : _GEN_760; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_762 = 6'h3a == cacheLine ? cache_58_line_0 : _GEN_761; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_763 = 6'h3b == cacheLine ? cache_59_line_0 : _GEN_762; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_764 = 6'h3c == cacheLine ? cache_60_line_0 : _GEN_763; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_765 = 6'h3d == cacheLine ? cache_61_line_0 : _GEN_764; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_766 = 6'h3e == cacheLine ? cache_62_line_0 : _GEN_765; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_767 = 6'h3f == cacheLine ? cache_63_line_0 : _GEN_766; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_769 = 6'h1 == cacheLine ? cache_1_line_3 : cache_0_line_3; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_770 = 6'h2 == cacheLine ? cache_2_line_3 : _GEN_769; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_771 = 6'h3 == cacheLine ? cache_3_line_3 : _GEN_770; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_772 = 6'h4 == cacheLine ? cache_4_line_3 : _GEN_771; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_773 = 6'h5 == cacheLine ? cache_5_line_3 : _GEN_772; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_774 = 6'h6 == cacheLine ? cache_6_line_3 : _GEN_773; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_775 = 6'h7 == cacheLine ? cache_7_line_3 : _GEN_774; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_776 = 6'h8 == cacheLine ? cache_8_line_3 : _GEN_775; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_777 = 6'h9 == cacheLine ? cache_9_line_3 : _GEN_776; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_778 = 6'ha == cacheLine ? cache_10_line_3 : _GEN_777; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_779 = 6'hb == cacheLine ? cache_11_line_3 : _GEN_778; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_780 = 6'hc == cacheLine ? cache_12_line_3 : _GEN_779; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_781 = 6'hd == cacheLine ? cache_13_line_3 : _GEN_780; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_782 = 6'he == cacheLine ? cache_14_line_3 : _GEN_781; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_783 = 6'hf == cacheLine ? cache_15_line_3 : _GEN_782; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_784 = 6'h10 == cacheLine ? cache_16_line_3 : _GEN_783; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_785 = 6'h11 == cacheLine ? cache_17_line_3 : _GEN_784; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_786 = 6'h12 == cacheLine ? cache_18_line_3 : _GEN_785; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_787 = 6'h13 == cacheLine ? cache_19_line_3 : _GEN_786; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_788 = 6'h14 == cacheLine ? cache_20_line_3 : _GEN_787; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_789 = 6'h15 == cacheLine ? cache_21_line_3 : _GEN_788; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_790 = 6'h16 == cacheLine ? cache_22_line_3 : _GEN_789; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_791 = 6'h17 == cacheLine ? cache_23_line_3 : _GEN_790; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_792 = 6'h18 == cacheLine ? cache_24_line_3 : _GEN_791; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_793 = 6'h19 == cacheLine ? cache_25_line_3 : _GEN_792; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_794 = 6'h1a == cacheLine ? cache_26_line_3 : _GEN_793; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_795 = 6'h1b == cacheLine ? cache_27_line_3 : _GEN_794; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_796 = 6'h1c == cacheLine ? cache_28_line_3 : _GEN_795; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_797 = 6'h1d == cacheLine ? cache_29_line_3 : _GEN_796; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_798 = 6'h1e == cacheLine ? cache_30_line_3 : _GEN_797; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_799 = 6'h1f == cacheLine ? cache_31_line_3 : _GEN_798; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_800 = 6'h20 == cacheLine ? cache_32_line_3 : _GEN_799; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_801 = 6'h21 == cacheLine ? cache_33_line_3 : _GEN_800; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_802 = 6'h22 == cacheLine ? cache_34_line_3 : _GEN_801; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_803 = 6'h23 == cacheLine ? cache_35_line_3 : _GEN_802; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_804 = 6'h24 == cacheLine ? cache_36_line_3 : _GEN_803; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_805 = 6'h25 == cacheLine ? cache_37_line_3 : _GEN_804; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_806 = 6'h26 == cacheLine ? cache_38_line_3 : _GEN_805; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_807 = 6'h27 == cacheLine ? cache_39_line_3 : _GEN_806; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_808 = 6'h28 == cacheLine ? cache_40_line_3 : _GEN_807; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_809 = 6'h29 == cacheLine ? cache_41_line_3 : _GEN_808; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_810 = 6'h2a == cacheLine ? cache_42_line_3 : _GEN_809; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_811 = 6'h2b == cacheLine ? cache_43_line_3 : _GEN_810; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_812 = 6'h2c == cacheLine ? cache_44_line_3 : _GEN_811; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_813 = 6'h2d == cacheLine ? cache_45_line_3 : _GEN_812; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_814 = 6'h2e == cacheLine ? cache_46_line_3 : _GEN_813; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_815 = 6'h2f == cacheLine ? cache_47_line_3 : _GEN_814; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_816 = 6'h30 == cacheLine ? cache_48_line_3 : _GEN_815; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_817 = 6'h31 == cacheLine ? cache_49_line_3 : _GEN_816; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_818 = 6'h32 == cacheLine ? cache_50_line_3 : _GEN_817; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_819 = 6'h33 == cacheLine ? cache_51_line_3 : _GEN_818; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_820 = 6'h34 == cacheLine ? cache_52_line_3 : _GEN_819; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_821 = 6'h35 == cacheLine ? cache_53_line_3 : _GEN_820; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_822 = 6'h36 == cacheLine ? cache_54_line_3 : _GEN_821; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_823 = 6'h37 == cacheLine ? cache_55_line_3 : _GEN_822; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_824 = 6'h38 == cacheLine ? cache_56_line_3 : _GEN_823; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_825 = 6'h39 == cacheLine ? cache_57_line_3 : _GEN_824; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_826 = 6'h3a == cacheLine ? cache_58_line_3 : _GEN_825; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_827 = 6'h3b == cacheLine ? cache_59_line_3 : _GEN_826; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_828 = 6'h3c == cacheLine ? cache_60_line_3 : _GEN_827; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_829 = 6'h3d == cacheLine ? cache_61_line_3 : _GEN_828; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_830 = 6'h3e == cacheLine ? cache_62_line_3 : _GEN_829; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_831 = 6'h3f == cacheLine ? cache_63_line_3 : _GEN_830; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_833 = 6'h1 == cacheLine ? cache_1_line_2 : cache_0_line_2; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_834 = 6'h2 == cacheLine ? cache_2_line_2 : _GEN_833; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_835 = 6'h3 == cacheLine ? cache_3_line_2 : _GEN_834; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_836 = 6'h4 == cacheLine ? cache_4_line_2 : _GEN_835; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_837 = 6'h5 == cacheLine ? cache_5_line_2 : _GEN_836; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_838 = 6'h6 == cacheLine ? cache_6_line_2 : _GEN_837; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_839 = 6'h7 == cacheLine ? cache_7_line_2 : _GEN_838; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_840 = 6'h8 == cacheLine ? cache_8_line_2 : _GEN_839; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_841 = 6'h9 == cacheLine ? cache_9_line_2 : _GEN_840; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_842 = 6'ha == cacheLine ? cache_10_line_2 : _GEN_841; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_843 = 6'hb == cacheLine ? cache_11_line_2 : _GEN_842; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_844 = 6'hc == cacheLine ? cache_12_line_2 : _GEN_843; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_845 = 6'hd == cacheLine ? cache_13_line_2 : _GEN_844; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_846 = 6'he == cacheLine ? cache_14_line_2 : _GEN_845; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_847 = 6'hf == cacheLine ? cache_15_line_2 : _GEN_846; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_848 = 6'h10 == cacheLine ? cache_16_line_2 : _GEN_847; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_849 = 6'h11 == cacheLine ? cache_17_line_2 : _GEN_848; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_850 = 6'h12 == cacheLine ? cache_18_line_2 : _GEN_849; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_851 = 6'h13 == cacheLine ? cache_19_line_2 : _GEN_850; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_852 = 6'h14 == cacheLine ? cache_20_line_2 : _GEN_851; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_853 = 6'h15 == cacheLine ? cache_21_line_2 : _GEN_852; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_854 = 6'h16 == cacheLine ? cache_22_line_2 : _GEN_853; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_855 = 6'h17 == cacheLine ? cache_23_line_2 : _GEN_854; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_856 = 6'h18 == cacheLine ? cache_24_line_2 : _GEN_855; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_857 = 6'h19 == cacheLine ? cache_25_line_2 : _GEN_856; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_858 = 6'h1a == cacheLine ? cache_26_line_2 : _GEN_857; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_859 = 6'h1b == cacheLine ? cache_27_line_2 : _GEN_858; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_860 = 6'h1c == cacheLine ? cache_28_line_2 : _GEN_859; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_861 = 6'h1d == cacheLine ? cache_29_line_2 : _GEN_860; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_862 = 6'h1e == cacheLine ? cache_30_line_2 : _GEN_861; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_863 = 6'h1f == cacheLine ? cache_31_line_2 : _GEN_862; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_864 = 6'h20 == cacheLine ? cache_32_line_2 : _GEN_863; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_865 = 6'h21 == cacheLine ? cache_33_line_2 : _GEN_864; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_866 = 6'h22 == cacheLine ? cache_34_line_2 : _GEN_865; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_867 = 6'h23 == cacheLine ? cache_35_line_2 : _GEN_866; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_868 = 6'h24 == cacheLine ? cache_36_line_2 : _GEN_867; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_869 = 6'h25 == cacheLine ? cache_37_line_2 : _GEN_868; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_870 = 6'h26 == cacheLine ? cache_38_line_2 : _GEN_869; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_871 = 6'h27 == cacheLine ? cache_39_line_2 : _GEN_870; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_872 = 6'h28 == cacheLine ? cache_40_line_2 : _GEN_871; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_873 = 6'h29 == cacheLine ? cache_41_line_2 : _GEN_872; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_874 = 6'h2a == cacheLine ? cache_42_line_2 : _GEN_873; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_875 = 6'h2b == cacheLine ? cache_43_line_2 : _GEN_874; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_876 = 6'h2c == cacheLine ? cache_44_line_2 : _GEN_875; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_877 = 6'h2d == cacheLine ? cache_45_line_2 : _GEN_876; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_878 = 6'h2e == cacheLine ? cache_46_line_2 : _GEN_877; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_879 = 6'h2f == cacheLine ? cache_47_line_2 : _GEN_878; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_880 = 6'h30 == cacheLine ? cache_48_line_2 : _GEN_879; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_881 = 6'h31 == cacheLine ? cache_49_line_2 : _GEN_880; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_882 = 6'h32 == cacheLine ? cache_50_line_2 : _GEN_881; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_883 = 6'h33 == cacheLine ? cache_51_line_2 : _GEN_882; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_884 = 6'h34 == cacheLine ? cache_52_line_2 : _GEN_883; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_885 = 6'h35 == cacheLine ? cache_53_line_2 : _GEN_884; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_886 = 6'h36 == cacheLine ? cache_54_line_2 : _GEN_885; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_887 = 6'h37 == cacheLine ? cache_55_line_2 : _GEN_886; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_888 = 6'h38 == cacheLine ? cache_56_line_2 : _GEN_887; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_889 = 6'h39 == cacheLine ? cache_57_line_2 : _GEN_888; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_890 = 6'h3a == cacheLine ? cache_58_line_2 : _GEN_889; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_891 = 6'h3b == cacheLine ? cache_59_line_2 : _GEN_890; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_892 = 6'h3c == cacheLine ? cache_60_line_2 : _GEN_891; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_893 = 6'h3d == cacheLine ? cache_61_line_2 : _GEN_892; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_894 = 6'h3e == cacheLine ? cache_62_line_2 : _GEN_893; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_895 = 6'h3f == cacheLine ? cache_63_line_2 : _GEN_894; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_897 = 6'h1 == cacheLine ? cache_1_line_5 : cache_0_line_5; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_898 = 6'h2 == cacheLine ? cache_2_line_5 : _GEN_897; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_899 = 6'h3 == cacheLine ? cache_3_line_5 : _GEN_898; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_900 = 6'h4 == cacheLine ? cache_4_line_5 : _GEN_899; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_901 = 6'h5 == cacheLine ? cache_5_line_5 : _GEN_900; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_902 = 6'h6 == cacheLine ? cache_6_line_5 : _GEN_901; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_903 = 6'h7 == cacheLine ? cache_7_line_5 : _GEN_902; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_904 = 6'h8 == cacheLine ? cache_8_line_5 : _GEN_903; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_905 = 6'h9 == cacheLine ? cache_9_line_5 : _GEN_904; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_906 = 6'ha == cacheLine ? cache_10_line_5 : _GEN_905; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_907 = 6'hb == cacheLine ? cache_11_line_5 : _GEN_906; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_908 = 6'hc == cacheLine ? cache_12_line_5 : _GEN_907; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_909 = 6'hd == cacheLine ? cache_13_line_5 : _GEN_908; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_910 = 6'he == cacheLine ? cache_14_line_5 : _GEN_909; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_911 = 6'hf == cacheLine ? cache_15_line_5 : _GEN_910; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_912 = 6'h10 == cacheLine ? cache_16_line_5 : _GEN_911; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_913 = 6'h11 == cacheLine ? cache_17_line_5 : _GEN_912; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_914 = 6'h12 == cacheLine ? cache_18_line_5 : _GEN_913; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_915 = 6'h13 == cacheLine ? cache_19_line_5 : _GEN_914; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_916 = 6'h14 == cacheLine ? cache_20_line_5 : _GEN_915; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_917 = 6'h15 == cacheLine ? cache_21_line_5 : _GEN_916; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_918 = 6'h16 == cacheLine ? cache_22_line_5 : _GEN_917; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_919 = 6'h17 == cacheLine ? cache_23_line_5 : _GEN_918; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_920 = 6'h18 == cacheLine ? cache_24_line_5 : _GEN_919; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_921 = 6'h19 == cacheLine ? cache_25_line_5 : _GEN_920; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_922 = 6'h1a == cacheLine ? cache_26_line_5 : _GEN_921; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_923 = 6'h1b == cacheLine ? cache_27_line_5 : _GEN_922; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_924 = 6'h1c == cacheLine ? cache_28_line_5 : _GEN_923; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_925 = 6'h1d == cacheLine ? cache_29_line_5 : _GEN_924; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_926 = 6'h1e == cacheLine ? cache_30_line_5 : _GEN_925; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_927 = 6'h1f == cacheLine ? cache_31_line_5 : _GEN_926; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_928 = 6'h20 == cacheLine ? cache_32_line_5 : _GEN_927; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_929 = 6'h21 == cacheLine ? cache_33_line_5 : _GEN_928; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_930 = 6'h22 == cacheLine ? cache_34_line_5 : _GEN_929; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_931 = 6'h23 == cacheLine ? cache_35_line_5 : _GEN_930; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_932 = 6'h24 == cacheLine ? cache_36_line_5 : _GEN_931; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_933 = 6'h25 == cacheLine ? cache_37_line_5 : _GEN_932; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_934 = 6'h26 == cacheLine ? cache_38_line_5 : _GEN_933; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_935 = 6'h27 == cacheLine ? cache_39_line_5 : _GEN_934; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_936 = 6'h28 == cacheLine ? cache_40_line_5 : _GEN_935; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_937 = 6'h29 == cacheLine ? cache_41_line_5 : _GEN_936; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_938 = 6'h2a == cacheLine ? cache_42_line_5 : _GEN_937; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_939 = 6'h2b == cacheLine ? cache_43_line_5 : _GEN_938; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_940 = 6'h2c == cacheLine ? cache_44_line_5 : _GEN_939; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_941 = 6'h2d == cacheLine ? cache_45_line_5 : _GEN_940; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_942 = 6'h2e == cacheLine ? cache_46_line_5 : _GEN_941; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_943 = 6'h2f == cacheLine ? cache_47_line_5 : _GEN_942; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_944 = 6'h30 == cacheLine ? cache_48_line_5 : _GEN_943; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_945 = 6'h31 == cacheLine ? cache_49_line_5 : _GEN_944; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_946 = 6'h32 == cacheLine ? cache_50_line_5 : _GEN_945; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_947 = 6'h33 == cacheLine ? cache_51_line_5 : _GEN_946; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_948 = 6'h34 == cacheLine ? cache_52_line_5 : _GEN_947; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_949 = 6'h35 == cacheLine ? cache_53_line_5 : _GEN_948; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_950 = 6'h36 == cacheLine ? cache_54_line_5 : _GEN_949; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_951 = 6'h37 == cacheLine ? cache_55_line_5 : _GEN_950; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_952 = 6'h38 == cacheLine ? cache_56_line_5 : _GEN_951; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_953 = 6'h39 == cacheLine ? cache_57_line_5 : _GEN_952; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_954 = 6'h3a == cacheLine ? cache_58_line_5 : _GEN_953; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_955 = 6'h3b == cacheLine ? cache_59_line_5 : _GEN_954; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_956 = 6'h3c == cacheLine ? cache_60_line_5 : _GEN_955; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_957 = 6'h3d == cacheLine ? cache_61_line_5 : _GEN_956; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_958 = 6'h3e == cacheLine ? cache_62_line_5 : _GEN_957; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_959 = 6'h3f == cacheLine ? cache_63_line_5 : _GEN_958; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_961 = 6'h1 == cacheLine ? cache_1_line_4 : cache_0_line_4; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_962 = 6'h2 == cacheLine ? cache_2_line_4 : _GEN_961; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_963 = 6'h3 == cacheLine ? cache_3_line_4 : _GEN_962; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_964 = 6'h4 == cacheLine ? cache_4_line_4 : _GEN_963; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_965 = 6'h5 == cacheLine ? cache_5_line_4 : _GEN_964; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_966 = 6'h6 == cacheLine ? cache_6_line_4 : _GEN_965; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_967 = 6'h7 == cacheLine ? cache_7_line_4 : _GEN_966; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_968 = 6'h8 == cacheLine ? cache_8_line_4 : _GEN_967; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_969 = 6'h9 == cacheLine ? cache_9_line_4 : _GEN_968; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_970 = 6'ha == cacheLine ? cache_10_line_4 : _GEN_969; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_971 = 6'hb == cacheLine ? cache_11_line_4 : _GEN_970; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_972 = 6'hc == cacheLine ? cache_12_line_4 : _GEN_971; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_973 = 6'hd == cacheLine ? cache_13_line_4 : _GEN_972; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_974 = 6'he == cacheLine ? cache_14_line_4 : _GEN_973; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_975 = 6'hf == cacheLine ? cache_15_line_4 : _GEN_974; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_976 = 6'h10 == cacheLine ? cache_16_line_4 : _GEN_975; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_977 = 6'h11 == cacheLine ? cache_17_line_4 : _GEN_976; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_978 = 6'h12 == cacheLine ? cache_18_line_4 : _GEN_977; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_979 = 6'h13 == cacheLine ? cache_19_line_4 : _GEN_978; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_980 = 6'h14 == cacheLine ? cache_20_line_4 : _GEN_979; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_981 = 6'h15 == cacheLine ? cache_21_line_4 : _GEN_980; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_982 = 6'h16 == cacheLine ? cache_22_line_4 : _GEN_981; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_983 = 6'h17 == cacheLine ? cache_23_line_4 : _GEN_982; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_984 = 6'h18 == cacheLine ? cache_24_line_4 : _GEN_983; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_985 = 6'h19 == cacheLine ? cache_25_line_4 : _GEN_984; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_986 = 6'h1a == cacheLine ? cache_26_line_4 : _GEN_985; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_987 = 6'h1b == cacheLine ? cache_27_line_4 : _GEN_986; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_988 = 6'h1c == cacheLine ? cache_28_line_4 : _GEN_987; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_989 = 6'h1d == cacheLine ? cache_29_line_4 : _GEN_988; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_990 = 6'h1e == cacheLine ? cache_30_line_4 : _GEN_989; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_991 = 6'h1f == cacheLine ? cache_31_line_4 : _GEN_990; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_992 = 6'h20 == cacheLine ? cache_32_line_4 : _GEN_991; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_993 = 6'h21 == cacheLine ? cache_33_line_4 : _GEN_992; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_994 = 6'h22 == cacheLine ? cache_34_line_4 : _GEN_993; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_995 = 6'h23 == cacheLine ? cache_35_line_4 : _GEN_994; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_996 = 6'h24 == cacheLine ? cache_36_line_4 : _GEN_995; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_997 = 6'h25 == cacheLine ? cache_37_line_4 : _GEN_996; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_998 = 6'h26 == cacheLine ? cache_38_line_4 : _GEN_997; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_999 = 6'h27 == cacheLine ? cache_39_line_4 : _GEN_998; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1000 = 6'h28 == cacheLine ? cache_40_line_4 : _GEN_999; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1001 = 6'h29 == cacheLine ? cache_41_line_4 : _GEN_1000; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1002 = 6'h2a == cacheLine ? cache_42_line_4 : _GEN_1001; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1003 = 6'h2b == cacheLine ? cache_43_line_4 : _GEN_1002; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1004 = 6'h2c == cacheLine ? cache_44_line_4 : _GEN_1003; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1005 = 6'h2d == cacheLine ? cache_45_line_4 : _GEN_1004; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1006 = 6'h2e == cacheLine ? cache_46_line_4 : _GEN_1005; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1007 = 6'h2f == cacheLine ? cache_47_line_4 : _GEN_1006; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1008 = 6'h30 == cacheLine ? cache_48_line_4 : _GEN_1007; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1009 = 6'h31 == cacheLine ? cache_49_line_4 : _GEN_1008; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1010 = 6'h32 == cacheLine ? cache_50_line_4 : _GEN_1009; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1011 = 6'h33 == cacheLine ? cache_51_line_4 : _GEN_1010; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1012 = 6'h34 == cacheLine ? cache_52_line_4 : _GEN_1011; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1013 = 6'h35 == cacheLine ? cache_53_line_4 : _GEN_1012; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1014 = 6'h36 == cacheLine ? cache_54_line_4 : _GEN_1013; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1015 = 6'h37 == cacheLine ? cache_55_line_4 : _GEN_1014; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1016 = 6'h38 == cacheLine ? cache_56_line_4 : _GEN_1015; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1017 = 6'h39 == cacheLine ? cache_57_line_4 : _GEN_1016; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1018 = 6'h3a == cacheLine ? cache_58_line_4 : _GEN_1017; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1019 = 6'h3b == cacheLine ? cache_59_line_4 : _GEN_1018; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1020 = 6'h3c == cacheLine ? cache_60_line_4 : _GEN_1019; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1021 = 6'h3d == cacheLine ? cache_61_line_4 : _GEN_1020; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1022 = 6'h3e == cacheLine ? cache_62_line_4 : _GEN_1021; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1023 = 6'h3f == cacheLine ? cache_63_line_4 : _GEN_1022; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1025 = 6'h1 == cacheLine ? cache_1_line_7 : cache_0_line_7; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1026 = 6'h2 == cacheLine ? cache_2_line_7 : _GEN_1025; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1027 = 6'h3 == cacheLine ? cache_3_line_7 : _GEN_1026; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1028 = 6'h4 == cacheLine ? cache_4_line_7 : _GEN_1027; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1029 = 6'h5 == cacheLine ? cache_5_line_7 : _GEN_1028; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1030 = 6'h6 == cacheLine ? cache_6_line_7 : _GEN_1029; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1031 = 6'h7 == cacheLine ? cache_7_line_7 : _GEN_1030; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1032 = 6'h8 == cacheLine ? cache_8_line_7 : _GEN_1031; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1033 = 6'h9 == cacheLine ? cache_9_line_7 : _GEN_1032; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1034 = 6'ha == cacheLine ? cache_10_line_7 : _GEN_1033; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1035 = 6'hb == cacheLine ? cache_11_line_7 : _GEN_1034; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1036 = 6'hc == cacheLine ? cache_12_line_7 : _GEN_1035; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1037 = 6'hd == cacheLine ? cache_13_line_7 : _GEN_1036; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1038 = 6'he == cacheLine ? cache_14_line_7 : _GEN_1037; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1039 = 6'hf == cacheLine ? cache_15_line_7 : _GEN_1038; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1040 = 6'h10 == cacheLine ? cache_16_line_7 : _GEN_1039; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1041 = 6'h11 == cacheLine ? cache_17_line_7 : _GEN_1040; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1042 = 6'h12 == cacheLine ? cache_18_line_7 : _GEN_1041; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1043 = 6'h13 == cacheLine ? cache_19_line_7 : _GEN_1042; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1044 = 6'h14 == cacheLine ? cache_20_line_7 : _GEN_1043; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1045 = 6'h15 == cacheLine ? cache_21_line_7 : _GEN_1044; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1046 = 6'h16 == cacheLine ? cache_22_line_7 : _GEN_1045; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1047 = 6'h17 == cacheLine ? cache_23_line_7 : _GEN_1046; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1048 = 6'h18 == cacheLine ? cache_24_line_7 : _GEN_1047; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1049 = 6'h19 == cacheLine ? cache_25_line_7 : _GEN_1048; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1050 = 6'h1a == cacheLine ? cache_26_line_7 : _GEN_1049; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1051 = 6'h1b == cacheLine ? cache_27_line_7 : _GEN_1050; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1052 = 6'h1c == cacheLine ? cache_28_line_7 : _GEN_1051; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1053 = 6'h1d == cacheLine ? cache_29_line_7 : _GEN_1052; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1054 = 6'h1e == cacheLine ? cache_30_line_7 : _GEN_1053; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1055 = 6'h1f == cacheLine ? cache_31_line_7 : _GEN_1054; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1056 = 6'h20 == cacheLine ? cache_32_line_7 : _GEN_1055; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1057 = 6'h21 == cacheLine ? cache_33_line_7 : _GEN_1056; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1058 = 6'h22 == cacheLine ? cache_34_line_7 : _GEN_1057; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1059 = 6'h23 == cacheLine ? cache_35_line_7 : _GEN_1058; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1060 = 6'h24 == cacheLine ? cache_36_line_7 : _GEN_1059; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1061 = 6'h25 == cacheLine ? cache_37_line_7 : _GEN_1060; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1062 = 6'h26 == cacheLine ? cache_38_line_7 : _GEN_1061; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1063 = 6'h27 == cacheLine ? cache_39_line_7 : _GEN_1062; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1064 = 6'h28 == cacheLine ? cache_40_line_7 : _GEN_1063; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1065 = 6'h29 == cacheLine ? cache_41_line_7 : _GEN_1064; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1066 = 6'h2a == cacheLine ? cache_42_line_7 : _GEN_1065; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1067 = 6'h2b == cacheLine ? cache_43_line_7 : _GEN_1066; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1068 = 6'h2c == cacheLine ? cache_44_line_7 : _GEN_1067; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1069 = 6'h2d == cacheLine ? cache_45_line_7 : _GEN_1068; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1070 = 6'h2e == cacheLine ? cache_46_line_7 : _GEN_1069; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1071 = 6'h2f == cacheLine ? cache_47_line_7 : _GEN_1070; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1072 = 6'h30 == cacheLine ? cache_48_line_7 : _GEN_1071; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1073 = 6'h31 == cacheLine ? cache_49_line_7 : _GEN_1072; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1074 = 6'h32 == cacheLine ? cache_50_line_7 : _GEN_1073; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1075 = 6'h33 == cacheLine ? cache_51_line_7 : _GEN_1074; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1076 = 6'h34 == cacheLine ? cache_52_line_7 : _GEN_1075; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1077 = 6'h35 == cacheLine ? cache_53_line_7 : _GEN_1076; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1078 = 6'h36 == cacheLine ? cache_54_line_7 : _GEN_1077; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1079 = 6'h37 == cacheLine ? cache_55_line_7 : _GEN_1078; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1080 = 6'h38 == cacheLine ? cache_56_line_7 : _GEN_1079; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1081 = 6'h39 == cacheLine ? cache_57_line_7 : _GEN_1080; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1082 = 6'h3a == cacheLine ? cache_58_line_7 : _GEN_1081; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1083 = 6'h3b == cacheLine ? cache_59_line_7 : _GEN_1082; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1084 = 6'h3c == cacheLine ? cache_60_line_7 : _GEN_1083; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1085 = 6'h3d == cacheLine ? cache_61_line_7 : _GEN_1084; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1086 = 6'h3e == cacheLine ? cache_62_line_7 : _GEN_1085; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1087 = 6'h3f == cacheLine ? cache_63_line_7 : _GEN_1086; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1089 = 6'h1 == cacheLine ? cache_1_line_6 : cache_0_line_6; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1090 = 6'h2 == cacheLine ? cache_2_line_6 : _GEN_1089; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1091 = 6'h3 == cacheLine ? cache_3_line_6 : _GEN_1090; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1092 = 6'h4 == cacheLine ? cache_4_line_6 : _GEN_1091; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1093 = 6'h5 == cacheLine ? cache_5_line_6 : _GEN_1092; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1094 = 6'h6 == cacheLine ? cache_6_line_6 : _GEN_1093; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1095 = 6'h7 == cacheLine ? cache_7_line_6 : _GEN_1094; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1096 = 6'h8 == cacheLine ? cache_8_line_6 : _GEN_1095; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1097 = 6'h9 == cacheLine ? cache_9_line_6 : _GEN_1096; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1098 = 6'ha == cacheLine ? cache_10_line_6 : _GEN_1097; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1099 = 6'hb == cacheLine ? cache_11_line_6 : _GEN_1098; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1100 = 6'hc == cacheLine ? cache_12_line_6 : _GEN_1099; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1101 = 6'hd == cacheLine ? cache_13_line_6 : _GEN_1100; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1102 = 6'he == cacheLine ? cache_14_line_6 : _GEN_1101; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1103 = 6'hf == cacheLine ? cache_15_line_6 : _GEN_1102; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1104 = 6'h10 == cacheLine ? cache_16_line_6 : _GEN_1103; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1105 = 6'h11 == cacheLine ? cache_17_line_6 : _GEN_1104; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1106 = 6'h12 == cacheLine ? cache_18_line_6 : _GEN_1105; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1107 = 6'h13 == cacheLine ? cache_19_line_6 : _GEN_1106; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1108 = 6'h14 == cacheLine ? cache_20_line_6 : _GEN_1107; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1109 = 6'h15 == cacheLine ? cache_21_line_6 : _GEN_1108; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1110 = 6'h16 == cacheLine ? cache_22_line_6 : _GEN_1109; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1111 = 6'h17 == cacheLine ? cache_23_line_6 : _GEN_1110; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1112 = 6'h18 == cacheLine ? cache_24_line_6 : _GEN_1111; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1113 = 6'h19 == cacheLine ? cache_25_line_6 : _GEN_1112; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1114 = 6'h1a == cacheLine ? cache_26_line_6 : _GEN_1113; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1115 = 6'h1b == cacheLine ? cache_27_line_6 : _GEN_1114; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1116 = 6'h1c == cacheLine ? cache_28_line_6 : _GEN_1115; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1117 = 6'h1d == cacheLine ? cache_29_line_6 : _GEN_1116; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1118 = 6'h1e == cacheLine ? cache_30_line_6 : _GEN_1117; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1119 = 6'h1f == cacheLine ? cache_31_line_6 : _GEN_1118; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1120 = 6'h20 == cacheLine ? cache_32_line_6 : _GEN_1119; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1121 = 6'h21 == cacheLine ? cache_33_line_6 : _GEN_1120; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1122 = 6'h22 == cacheLine ? cache_34_line_6 : _GEN_1121; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1123 = 6'h23 == cacheLine ? cache_35_line_6 : _GEN_1122; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1124 = 6'h24 == cacheLine ? cache_36_line_6 : _GEN_1123; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1125 = 6'h25 == cacheLine ? cache_37_line_6 : _GEN_1124; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1126 = 6'h26 == cacheLine ? cache_38_line_6 : _GEN_1125; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1127 = 6'h27 == cacheLine ? cache_39_line_6 : _GEN_1126; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1128 = 6'h28 == cacheLine ? cache_40_line_6 : _GEN_1127; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1129 = 6'h29 == cacheLine ? cache_41_line_6 : _GEN_1128; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1130 = 6'h2a == cacheLine ? cache_42_line_6 : _GEN_1129; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1131 = 6'h2b == cacheLine ? cache_43_line_6 : _GEN_1130; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1132 = 6'h2c == cacheLine ? cache_44_line_6 : _GEN_1131; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1133 = 6'h2d == cacheLine ? cache_45_line_6 : _GEN_1132; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1134 = 6'h2e == cacheLine ? cache_46_line_6 : _GEN_1133; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1135 = 6'h2f == cacheLine ? cache_47_line_6 : _GEN_1134; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1136 = 6'h30 == cacheLine ? cache_48_line_6 : _GEN_1135; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1137 = 6'h31 == cacheLine ? cache_49_line_6 : _GEN_1136; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1138 = 6'h32 == cacheLine ? cache_50_line_6 : _GEN_1137; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1139 = 6'h33 == cacheLine ? cache_51_line_6 : _GEN_1138; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1140 = 6'h34 == cacheLine ? cache_52_line_6 : _GEN_1139; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1141 = 6'h35 == cacheLine ? cache_53_line_6 : _GEN_1140; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1142 = 6'h36 == cacheLine ? cache_54_line_6 : _GEN_1141; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1143 = 6'h37 == cacheLine ? cache_55_line_6 : _GEN_1142; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1144 = 6'h38 == cacheLine ? cache_56_line_6 : _GEN_1143; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1145 = 6'h39 == cacheLine ? cache_57_line_6 : _GEN_1144; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1146 = 6'h3a == cacheLine ? cache_58_line_6 : _GEN_1145; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1147 = 6'h3b == cacheLine ? cache_59_line_6 : _GEN_1146; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1148 = 6'h3c == cacheLine ? cache_60_line_6 : _GEN_1147; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1149 = 6'h3d == cacheLine ? cache_61_line_6 : _GEN_1148; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1150 = 6'h3e == cacheLine ? cache_62_line_6 : _GEN_1149; // @[Cache.scala 45:{39,39}]
  wire [31:0] _GEN_1151 = 6'h3f == cacheLine ? cache_63_line_6 : _GEN_1150; // @[Cache.scala 45:{39,39}]
  wire [255:0] _dataBuffer_T = {_GEN_1087,_GEN_1151,_GEN_959,_GEN_1023,_GEN_831,_GEN_895,_GEN_703,_GEN_767}; // @[Cache.scala 45:39]
  wire  _GEN_1152 = _GEN_3972 | cache_0_validBit; // @[Cache.scala 32:22 49:{31,31}]
  wire  _GEN_1153 = _GEN_3986 | cache_1_validBit; // @[Cache.scala 32:22 49:{31,31}]
  wire  _GEN_1154 = _GEN_4002 | cache_2_validBit; // @[Cache.scala 32:22 49:{31,31}]
  wire  _GEN_1155 = _GEN_4018 | cache_3_validBit; // @[Cache.scala 32:22 49:{31,31}]
  wire  _GEN_1156 = _GEN_4034 | cache_4_validBit; // @[Cache.scala 32:22 49:{31,31}]
  wire  _GEN_1157 = _GEN_4050 | cache_5_validBit; // @[Cache.scala 32:22 49:{31,31}]
  wire  _GEN_1158 = _GEN_4066 | cache_6_validBit; // @[Cache.scala 32:22 49:{31,31}]
  wire  _GEN_1159 = _GEN_4082 | cache_7_validBit; // @[Cache.scala 32:22 49:{31,31}]
  wire  _GEN_1160 = _GEN_4098 | cache_8_validBit; // @[Cache.scala 32:22 49:{31,31}]
  wire  _GEN_1161 = _GEN_4114 | cache_9_validBit; // @[Cache.scala 32:22 49:{31,31}]
  wire  _GEN_1162 = _GEN_4130 | cache_10_validBit; // @[Cache.scala 32:22 49:{31,31}]
  wire  _GEN_1163 = _GEN_4146 | cache_11_validBit; // @[Cache.scala 32:22 49:{31,31}]
  wire  _GEN_1164 = _GEN_4162 | cache_12_validBit; // @[Cache.scala 32:22 49:{31,31}]
  wire  _GEN_1165 = _GEN_4178 | cache_13_validBit; // @[Cache.scala 32:22 49:{31,31}]
  wire  _GEN_1166 = _GEN_4194 | cache_14_validBit; // @[Cache.scala 32:22 49:{31,31}]
  wire  _GEN_1167 = _GEN_4210 | cache_15_validBit; // @[Cache.scala 32:22 49:{31,31}]
  wire  _GEN_1168 = _GEN_4226 | cache_16_validBit; // @[Cache.scala 32:22 49:{31,31}]
  wire  _GEN_1169 = _GEN_4242 | cache_17_validBit; // @[Cache.scala 32:22 49:{31,31}]
  wire  _GEN_1170 = _GEN_4258 | cache_18_validBit; // @[Cache.scala 32:22 49:{31,31}]
  wire  _GEN_1171 = _GEN_4274 | cache_19_validBit; // @[Cache.scala 32:22 49:{31,31}]
  wire  _GEN_1172 = _GEN_4290 | cache_20_validBit; // @[Cache.scala 32:22 49:{31,31}]
  wire  _GEN_1173 = _GEN_4306 | cache_21_validBit; // @[Cache.scala 32:22 49:{31,31}]
  wire  _GEN_1174 = _GEN_4322 | cache_22_validBit; // @[Cache.scala 32:22 49:{31,31}]
  wire  _GEN_1175 = _GEN_4338 | cache_23_validBit; // @[Cache.scala 32:22 49:{31,31}]
  wire  _GEN_1176 = _GEN_4354 | cache_24_validBit; // @[Cache.scala 32:22 49:{31,31}]
  wire  _GEN_1177 = _GEN_4370 | cache_25_validBit; // @[Cache.scala 32:22 49:{31,31}]
  wire  _GEN_1178 = _GEN_4386 | cache_26_validBit; // @[Cache.scala 32:22 49:{31,31}]
  wire  _GEN_1179 = _GEN_4402 | cache_27_validBit; // @[Cache.scala 32:22 49:{31,31}]
  wire  _GEN_1180 = _GEN_4418 | cache_28_validBit; // @[Cache.scala 32:22 49:{31,31}]
  wire  _GEN_1181 = _GEN_4434 | cache_29_validBit; // @[Cache.scala 32:22 49:{31,31}]
  wire  _GEN_1182 = _GEN_4450 | cache_30_validBit; // @[Cache.scala 32:22 49:{31,31}]
  wire  _GEN_1183 = _GEN_4466 | cache_31_validBit; // @[Cache.scala 32:22 49:{31,31}]
  wire  _GEN_1184 = _GEN_4482 | cache_32_validBit; // @[Cache.scala 32:22 49:{31,31}]
  wire  _GEN_1185 = _GEN_4498 | cache_33_validBit; // @[Cache.scala 32:22 49:{31,31}]
  wire  _GEN_1186 = _GEN_4514 | cache_34_validBit; // @[Cache.scala 32:22 49:{31,31}]
  wire  _GEN_1187 = _GEN_4530 | cache_35_validBit; // @[Cache.scala 32:22 49:{31,31}]
  wire  _GEN_1188 = _GEN_4546 | cache_36_validBit; // @[Cache.scala 32:22 49:{31,31}]
  wire  _GEN_1189 = _GEN_4562 | cache_37_validBit; // @[Cache.scala 32:22 49:{31,31}]
  wire  _GEN_1190 = _GEN_4578 | cache_38_validBit; // @[Cache.scala 32:22 49:{31,31}]
  wire  _GEN_1191 = _GEN_4594 | cache_39_validBit; // @[Cache.scala 32:22 49:{31,31}]
  wire  _GEN_1192 = _GEN_4610 | cache_40_validBit; // @[Cache.scala 32:22 49:{31,31}]
  wire  _GEN_1193 = _GEN_4626 | cache_41_validBit; // @[Cache.scala 32:22 49:{31,31}]
  wire  _GEN_1194 = _GEN_4642 | cache_42_validBit; // @[Cache.scala 32:22 49:{31,31}]
  wire  _GEN_1195 = _GEN_4658 | cache_43_validBit; // @[Cache.scala 32:22 49:{31,31}]
  wire  _GEN_1196 = _GEN_4674 | cache_44_validBit; // @[Cache.scala 32:22 49:{31,31}]
  wire  _GEN_1197 = _GEN_4690 | cache_45_validBit; // @[Cache.scala 32:22 49:{31,31}]
  wire  _GEN_1198 = _GEN_4706 | cache_46_validBit; // @[Cache.scala 32:22 49:{31,31}]
  wire  _GEN_1199 = _GEN_4722 | cache_47_validBit; // @[Cache.scala 32:22 49:{31,31}]
  wire  _GEN_1200 = _GEN_4738 | cache_48_validBit; // @[Cache.scala 32:22 49:{31,31}]
  wire  _GEN_1201 = _GEN_4754 | cache_49_validBit; // @[Cache.scala 32:22 49:{31,31}]
  wire  _GEN_1202 = _GEN_4770 | cache_50_validBit; // @[Cache.scala 32:22 49:{31,31}]
  wire  _GEN_1203 = _GEN_4786 | cache_51_validBit; // @[Cache.scala 32:22 49:{31,31}]
  wire  _GEN_1204 = _GEN_4802 | cache_52_validBit; // @[Cache.scala 32:22 49:{31,31}]
  wire  _GEN_1205 = _GEN_4818 | cache_53_validBit; // @[Cache.scala 32:22 49:{31,31}]
  wire  _GEN_1206 = _GEN_4834 | cache_54_validBit; // @[Cache.scala 32:22 49:{31,31}]
  wire  _GEN_1207 = _GEN_4850 | cache_55_validBit; // @[Cache.scala 32:22 49:{31,31}]
  wire  _GEN_1208 = _GEN_4866 | cache_56_validBit; // @[Cache.scala 32:22 49:{31,31}]
  wire  _GEN_1209 = _GEN_4882 | cache_57_validBit; // @[Cache.scala 32:22 49:{31,31}]
  wire  _GEN_1210 = _GEN_4898 | cache_58_validBit; // @[Cache.scala 32:22 49:{31,31}]
  wire  _GEN_1211 = _GEN_4914 | cache_59_validBit; // @[Cache.scala 32:22 49:{31,31}]
  wire  _GEN_1212 = _GEN_4930 | cache_60_validBit; // @[Cache.scala 32:22 49:{31,31}]
  wire  _GEN_1213 = _GEN_4946 | cache_61_validBit; // @[Cache.scala 32:22 49:{31,31}]
  wire  _GEN_1214 = _GEN_4962 | cache_62_validBit; // @[Cache.scala 32:22 49:{31,31}]
  wire  _GEN_1215 = _GEN_4978 | cache_63_validBit; // @[Cache.scala 32:22 49:{31,31}]
  wire [31:0] _GEN_1280 = 6'h0 == cacheLine ? io_writeBlock[31:0] : cache_0_line_0; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1281 = 6'h1 == cacheLine ? io_writeBlock[31:0] : cache_1_line_0; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1282 = 6'h2 == cacheLine ? io_writeBlock[31:0] : cache_2_line_0; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1283 = 6'h3 == cacheLine ? io_writeBlock[31:0] : cache_3_line_0; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1284 = 6'h4 == cacheLine ? io_writeBlock[31:0] : cache_4_line_0; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1285 = 6'h5 == cacheLine ? io_writeBlock[31:0] : cache_5_line_0; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1286 = 6'h6 == cacheLine ? io_writeBlock[31:0] : cache_6_line_0; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1287 = 6'h7 == cacheLine ? io_writeBlock[31:0] : cache_7_line_0; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1288 = 6'h8 == cacheLine ? io_writeBlock[31:0] : cache_8_line_0; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1289 = 6'h9 == cacheLine ? io_writeBlock[31:0] : cache_9_line_0; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1290 = 6'ha == cacheLine ? io_writeBlock[31:0] : cache_10_line_0; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1291 = 6'hb == cacheLine ? io_writeBlock[31:0] : cache_11_line_0; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1292 = 6'hc == cacheLine ? io_writeBlock[31:0] : cache_12_line_0; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1293 = 6'hd == cacheLine ? io_writeBlock[31:0] : cache_13_line_0; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1294 = 6'he == cacheLine ? io_writeBlock[31:0] : cache_14_line_0; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1295 = 6'hf == cacheLine ? io_writeBlock[31:0] : cache_15_line_0; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1296 = 6'h10 == cacheLine ? io_writeBlock[31:0] : cache_16_line_0; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1297 = 6'h11 == cacheLine ? io_writeBlock[31:0] : cache_17_line_0; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1298 = 6'h12 == cacheLine ? io_writeBlock[31:0] : cache_18_line_0; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1299 = 6'h13 == cacheLine ? io_writeBlock[31:0] : cache_19_line_0; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1300 = 6'h14 == cacheLine ? io_writeBlock[31:0] : cache_20_line_0; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1301 = 6'h15 == cacheLine ? io_writeBlock[31:0] : cache_21_line_0; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1302 = 6'h16 == cacheLine ? io_writeBlock[31:0] : cache_22_line_0; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1303 = 6'h17 == cacheLine ? io_writeBlock[31:0] : cache_23_line_0; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1304 = 6'h18 == cacheLine ? io_writeBlock[31:0] : cache_24_line_0; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1305 = 6'h19 == cacheLine ? io_writeBlock[31:0] : cache_25_line_0; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1306 = 6'h1a == cacheLine ? io_writeBlock[31:0] : cache_26_line_0; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1307 = 6'h1b == cacheLine ? io_writeBlock[31:0] : cache_27_line_0; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1308 = 6'h1c == cacheLine ? io_writeBlock[31:0] : cache_28_line_0; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1309 = 6'h1d == cacheLine ? io_writeBlock[31:0] : cache_29_line_0; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1310 = 6'h1e == cacheLine ? io_writeBlock[31:0] : cache_30_line_0; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1311 = 6'h1f == cacheLine ? io_writeBlock[31:0] : cache_31_line_0; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1312 = 6'h20 == cacheLine ? io_writeBlock[31:0] : cache_32_line_0; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1313 = 6'h21 == cacheLine ? io_writeBlock[31:0] : cache_33_line_0; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1314 = 6'h22 == cacheLine ? io_writeBlock[31:0] : cache_34_line_0; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1315 = 6'h23 == cacheLine ? io_writeBlock[31:0] : cache_35_line_0; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1316 = 6'h24 == cacheLine ? io_writeBlock[31:0] : cache_36_line_0; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1317 = 6'h25 == cacheLine ? io_writeBlock[31:0] : cache_37_line_0; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1318 = 6'h26 == cacheLine ? io_writeBlock[31:0] : cache_38_line_0; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1319 = 6'h27 == cacheLine ? io_writeBlock[31:0] : cache_39_line_0; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1320 = 6'h28 == cacheLine ? io_writeBlock[31:0] : cache_40_line_0; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1321 = 6'h29 == cacheLine ? io_writeBlock[31:0] : cache_41_line_0; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1322 = 6'h2a == cacheLine ? io_writeBlock[31:0] : cache_42_line_0; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1323 = 6'h2b == cacheLine ? io_writeBlock[31:0] : cache_43_line_0; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1324 = 6'h2c == cacheLine ? io_writeBlock[31:0] : cache_44_line_0; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1325 = 6'h2d == cacheLine ? io_writeBlock[31:0] : cache_45_line_0; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1326 = 6'h2e == cacheLine ? io_writeBlock[31:0] : cache_46_line_0; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1327 = 6'h2f == cacheLine ? io_writeBlock[31:0] : cache_47_line_0; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1328 = 6'h30 == cacheLine ? io_writeBlock[31:0] : cache_48_line_0; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1329 = 6'h31 == cacheLine ? io_writeBlock[31:0] : cache_49_line_0; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1330 = 6'h32 == cacheLine ? io_writeBlock[31:0] : cache_50_line_0; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1331 = 6'h33 == cacheLine ? io_writeBlock[31:0] : cache_51_line_0; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1332 = 6'h34 == cacheLine ? io_writeBlock[31:0] : cache_52_line_0; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1333 = 6'h35 == cacheLine ? io_writeBlock[31:0] : cache_53_line_0; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1334 = 6'h36 == cacheLine ? io_writeBlock[31:0] : cache_54_line_0; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1335 = 6'h37 == cacheLine ? io_writeBlock[31:0] : cache_55_line_0; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1336 = 6'h38 == cacheLine ? io_writeBlock[31:0] : cache_56_line_0; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1337 = 6'h39 == cacheLine ? io_writeBlock[31:0] : cache_57_line_0; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1338 = 6'h3a == cacheLine ? io_writeBlock[31:0] : cache_58_line_0; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1339 = 6'h3b == cacheLine ? io_writeBlock[31:0] : cache_59_line_0; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1340 = 6'h3c == cacheLine ? io_writeBlock[31:0] : cache_60_line_0; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1341 = 6'h3d == cacheLine ? io_writeBlock[31:0] : cache_61_line_0; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1342 = 6'h3e == cacheLine ? io_writeBlock[31:0] : cache_62_line_0; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1343 = 6'h3f == cacheLine ? io_writeBlock[31:0] : cache_63_line_0; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1344 = 6'h0 == cacheLine ? io_writeBlock[63:32] : cache_0_line_1; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1345 = 6'h1 == cacheLine ? io_writeBlock[63:32] : cache_1_line_1; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1346 = 6'h2 == cacheLine ? io_writeBlock[63:32] : cache_2_line_1; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1347 = 6'h3 == cacheLine ? io_writeBlock[63:32] : cache_3_line_1; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1348 = 6'h4 == cacheLine ? io_writeBlock[63:32] : cache_4_line_1; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1349 = 6'h5 == cacheLine ? io_writeBlock[63:32] : cache_5_line_1; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1350 = 6'h6 == cacheLine ? io_writeBlock[63:32] : cache_6_line_1; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1351 = 6'h7 == cacheLine ? io_writeBlock[63:32] : cache_7_line_1; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1352 = 6'h8 == cacheLine ? io_writeBlock[63:32] : cache_8_line_1; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1353 = 6'h9 == cacheLine ? io_writeBlock[63:32] : cache_9_line_1; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1354 = 6'ha == cacheLine ? io_writeBlock[63:32] : cache_10_line_1; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1355 = 6'hb == cacheLine ? io_writeBlock[63:32] : cache_11_line_1; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1356 = 6'hc == cacheLine ? io_writeBlock[63:32] : cache_12_line_1; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1357 = 6'hd == cacheLine ? io_writeBlock[63:32] : cache_13_line_1; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1358 = 6'he == cacheLine ? io_writeBlock[63:32] : cache_14_line_1; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1359 = 6'hf == cacheLine ? io_writeBlock[63:32] : cache_15_line_1; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1360 = 6'h10 == cacheLine ? io_writeBlock[63:32] : cache_16_line_1; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1361 = 6'h11 == cacheLine ? io_writeBlock[63:32] : cache_17_line_1; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1362 = 6'h12 == cacheLine ? io_writeBlock[63:32] : cache_18_line_1; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1363 = 6'h13 == cacheLine ? io_writeBlock[63:32] : cache_19_line_1; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1364 = 6'h14 == cacheLine ? io_writeBlock[63:32] : cache_20_line_1; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1365 = 6'h15 == cacheLine ? io_writeBlock[63:32] : cache_21_line_1; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1366 = 6'h16 == cacheLine ? io_writeBlock[63:32] : cache_22_line_1; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1367 = 6'h17 == cacheLine ? io_writeBlock[63:32] : cache_23_line_1; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1368 = 6'h18 == cacheLine ? io_writeBlock[63:32] : cache_24_line_1; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1369 = 6'h19 == cacheLine ? io_writeBlock[63:32] : cache_25_line_1; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1370 = 6'h1a == cacheLine ? io_writeBlock[63:32] : cache_26_line_1; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1371 = 6'h1b == cacheLine ? io_writeBlock[63:32] : cache_27_line_1; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1372 = 6'h1c == cacheLine ? io_writeBlock[63:32] : cache_28_line_1; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1373 = 6'h1d == cacheLine ? io_writeBlock[63:32] : cache_29_line_1; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1374 = 6'h1e == cacheLine ? io_writeBlock[63:32] : cache_30_line_1; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1375 = 6'h1f == cacheLine ? io_writeBlock[63:32] : cache_31_line_1; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1376 = 6'h20 == cacheLine ? io_writeBlock[63:32] : cache_32_line_1; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1377 = 6'h21 == cacheLine ? io_writeBlock[63:32] : cache_33_line_1; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1378 = 6'h22 == cacheLine ? io_writeBlock[63:32] : cache_34_line_1; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1379 = 6'h23 == cacheLine ? io_writeBlock[63:32] : cache_35_line_1; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1380 = 6'h24 == cacheLine ? io_writeBlock[63:32] : cache_36_line_1; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1381 = 6'h25 == cacheLine ? io_writeBlock[63:32] : cache_37_line_1; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1382 = 6'h26 == cacheLine ? io_writeBlock[63:32] : cache_38_line_1; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1383 = 6'h27 == cacheLine ? io_writeBlock[63:32] : cache_39_line_1; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1384 = 6'h28 == cacheLine ? io_writeBlock[63:32] : cache_40_line_1; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1385 = 6'h29 == cacheLine ? io_writeBlock[63:32] : cache_41_line_1; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1386 = 6'h2a == cacheLine ? io_writeBlock[63:32] : cache_42_line_1; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1387 = 6'h2b == cacheLine ? io_writeBlock[63:32] : cache_43_line_1; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1388 = 6'h2c == cacheLine ? io_writeBlock[63:32] : cache_44_line_1; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1389 = 6'h2d == cacheLine ? io_writeBlock[63:32] : cache_45_line_1; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1390 = 6'h2e == cacheLine ? io_writeBlock[63:32] : cache_46_line_1; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1391 = 6'h2f == cacheLine ? io_writeBlock[63:32] : cache_47_line_1; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1392 = 6'h30 == cacheLine ? io_writeBlock[63:32] : cache_48_line_1; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1393 = 6'h31 == cacheLine ? io_writeBlock[63:32] : cache_49_line_1; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1394 = 6'h32 == cacheLine ? io_writeBlock[63:32] : cache_50_line_1; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1395 = 6'h33 == cacheLine ? io_writeBlock[63:32] : cache_51_line_1; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1396 = 6'h34 == cacheLine ? io_writeBlock[63:32] : cache_52_line_1; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1397 = 6'h35 == cacheLine ? io_writeBlock[63:32] : cache_53_line_1; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1398 = 6'h36 == cacheLine ? io_writeBlock[63:32] : cache_54_line_1; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1399 = 6'h37 == cacheLine ? io_writeBlock[63:32] : cache_55_line_1; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1400 = 6'h38 == cacheLine ? io_writeBlock[63:32] : cache_56_line_1; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1401 = 6'h39 == cacheLine ? io_writeBlock[63:32] : cache_57_line_1; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1402 = 6'h3a == cacheLine ? io_writeBlock[63:32] : cache_58_line_1; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1403 = 6'h3b == cacheLine ? io_writeBlock[63:32] : cache_59_line_1; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1404 = 6'h3c == cacheLine ? io_writeBlock[63:32] : cache_60_line_1; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1405 = 6'h3d == cacheLine ? io_writeBlock[63:32] : cache_61_line_1; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1406 = 6'h3e == cacheLine ? io_writeBlock[63:32] : cache_62_line_1; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1407 = 6'h3f == cacheLine ? io_writeBlock[63:32] : cache_63_line_1; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1408 = 6'h0 == cacheLine ? io_writeBlock[95:64] : cache_0_line_2; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1409 = 6'h1 == cacheLine ? io_writeBlock[95:64] : cache_1_line_2; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1410 = 6'h2 == cacheLine ? io_writeBlock[95:64] : cache_2_line_2; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1411 = 6'h3 == cacheLine ? io_writeBlock[95:64] : cache_3_line_2; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1412 = 6'h4 == cacheLine ? io_writeBlock[95:64] : cache_4_line_2; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1413 = 6'h5 == cacheLine ? io_writeBlock[95:64] : cache_5_line_2; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1414 = 6'h6 == cacheLine ? io_writeBlock[95:64] : cache_6_line_2; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1415 = 6'h7 == cacheLine ? io_writeBlock[95:64] : cache_7_line_2; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1416 = 6'h8 == cacheLine ? io_writeBlock[95:64] : cache_8_line_2; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1417 = 6'h9 == cacheLine ? io_writeBlock[95:64] : cache_9_line_2; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1418 = 6'ha == cacheLine ? io_writeBlock[95:64] : cache_10_line_2; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1419 = 6'hb == cacheLine ? io_writeBlock[95:64] : cache_11_line_2; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1420 = 6'hc == cacheLine ? io_writeBlock[95:64] : cache_12_line_2; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1421 = 6'hd == cacheLine ? io_writeBlock[95:64] : cache_13_line_2; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1422 = 6'he == cacheLine ? io_writeBlock[95:64] : cache_14_line_2; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1423 = 6'hf == cacheLine ? io_writeBlock[95:64] : cache_15_line_2; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1424 = 6'h10 == cacheLine ? io_writeBlock[95:64] : cache_16_line_2; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1425 = 6'h11 == cacheLine ? io_writeBlock[95:64] : cache_17_line_2; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1426 = 6'h12 == cacheLine ? io_writeBlock[95:64] : cache_18_line_2; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1427 = 6'h13 == cacheLine ? io_writeBlock[95:64] : cache_19_line_2; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1428 = 6'h14 == cacheLine ? io_writeBlock[95:64] : cache_20_line_2; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1429 = 6'h15 == cacheLine ? io_writeBlock[95:64] : cache_21_line_2; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1430 = 6'h16 == cacheLine ? io_writeBlock[95:64] : cache_22_line_2; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1431 = 6'h17 == cacheLine ? io_writeBlock[95:64] : cache_23_line_2; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1432 = 6'h18 == cacheLine ? io_writeBlock[95:64] : cache_24_line_2; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1433 = 6'h19 == cacheLine ? io_writeBlock[95:64] : cache_25_line_2; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1434 = 6'h1a == cacheLine ? io_writeBlock[95:64] : cache_26_line_2; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1435 = 6'h1b == cacheLine ? io_writeBlock[95:64] : cache_27_line_2; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1436 = 6'h1c == cacheLine ? io_writeBlock[95:64] : cache_28_line_2; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1437 = 6'h1d == cacheLine ? io_writeBlock[95:64] : cache_29_line_2; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1438 = 6'h1e == cacheLine ? io_writeBlock[95:64] : cache_30_line_2; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1439 = 6'h1f == cacheLine ? io_writeBlock[95:64] : cache_31_line_2; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1440 = 6'h20 == cacheLine ? io_writeBlock[95:64] : cache_32_line_2; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1441 = 6'h21 == cacheLine ? io_writeBlock[95:64] : cache_33_line_2; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1442 = 6'h22 == cacheLine ? io_writeBlock[95:64] : cache_34_line_2; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1443 = 6'h23 == cacheLine ? io_writeBlock[95:64] : cache_35_line_2; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1444 = 6'h24 == cacheLine ? io_writeBlock[95:64] : cache_36_line_2; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1445 = 6'h25 == cacheLine ? io_writeBlock[95:64] : cache_37_line_2; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1446 = 6'h26 == cacheLine ? io_writeBlock[95:64] : cache_38_line_2; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1447 = 6'h27 == cacheLine ? io_writeBlock[95:64] : cache_39_line_2; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1448 = 6'h28 == cacheLine ? io_writeBlock[95:64] : cache_40_line_2; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1449 = 6'h29 == cacheLine ? io_writeBlock[95:64] : cache_41_line_2; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1450 = 6'h2a == cacheLine ? io_writeBlock[95:64] : cache_42_line_2; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1451 = 6'h2b == cacheLine ? io_writeBlock[95:64] : cache_43_line_2; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1452 = 6'h2c == cacheLine ? io_writeBlock[95:64] : cache_44_line_2; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1453 = 6'h2d == cacheLine ? io_writeBlock[95:64] : cache_45_line_2; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1454 = 6'h2e == cacheLine ? io_writeBlock[95:64] : cache_46_line_2; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1455 = 6'h2f == cacheLine ? io_writeBlock[95:64] : cache_47_line_2; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1456 = 6'h30 == cacheLine ? io_writeBlock[95:64] : cache_48_line_2; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1457 = 6'h31 == cacheLine ? io_writeBlock[95:64] : cache_49_line_2; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1458 = 6'h32 == cacheLine ? io_writeBlock[95:64] : cache_50_line_2; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1459 = 6'h33 == cacheLine ? io_writeBlock[95:64] : cache_51_line_2; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1460 = 6'h34 == cacheLine ? io_writeBlock[95:64] : cache_52_line_2; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1461 = 6'h35 == cacheLine ? io_writeBlock[95:64] : cache_53_line_2; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1462 = 6'h36 == cacheLine ? io_writeBlock[95:64] : cache_54_line_2; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1463 = 6'h37 == cacheLine ? io_writeBlock[95:64] : cache_55_line_2; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1464 = 6'h38 == cacheLine ? io_writeBlock[95:64] : cache_56_line_2; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1465 = 6'h39 == cacheLine ? io_writeBlock[95:64] : cache_57_line_2; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1466 = 6'h3a == cacheLine ? io_writeBlock[95:64] : cache_58_line_2; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1467 = 6'h3b == cacheLine ? io_writeBlock[95:64] : cache_59_line_2; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1468 = 6'h3c == cacheLine ? io_writeBlock[95:64] : cache_60_line_2; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1469 = 6'h3d == cacheLine ? io_writeBlock[95:64] : cache_61_line_2; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1470 = 6'h3e == cacheLine ? io_writeBlock[95:64] : cache_62_line_2; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1471 = 6'h3f == cacheLine ? io_writeBlock[95:64] : cache_63_line_2; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1472 = 6'h0 == cacheLine ? io_writeBlock[127:96] : cache_0_line_3; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1473 = 6'h1 == cacheLine ? io_writeBlock[127:96] : cache_1_line_3; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1474 = 6'h2 == cacheLine ? io_writeBlock[127:96] : cache_2_line_3; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1475 = 6'h3 == cacheLine ? io_writeBlock[127:96] : cache_3_line_3; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1476 = 6'h4 == cacheLine ? io_writeBlock[127:96] : cache_4_line_3; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1477 = 6'h5 == cacheLine ? io_writeBlock[127:96] : cache_5_line_3; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1478 = 6'h6 == cacheLine ? io_writeBlock[127:96] : cache_6_line_3; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1479 = 6'h7 == cacheLine ? io_writeBlock[127:96] : cache_7_line_3; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1480 = 6'h8 == cacheLine ? io_writeBlock[127:96] : cache_8_line_3; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1481 = 6'h9 == cacheLine ? io_writeBlock[127:96] : cache_9_line_3; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1482 = 6'ha == cacheLine ? io_writeBlock[127:96] : cache_10_line_3; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1483 = 6'hb == cacheLine ? io_writeBlock[127:96] : cache_11_line_3; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1484 = 6'hc == cacheLine ? io_writeBlock[127:96] : cache_12_line_3; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1485 = 6'hd == cacheLine ? io_writeBlock[127:96] : cache_13_line_3; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1486 = 6'he == cacheLine ? io_writeBlock[127:96] : cache_14_line_3; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1487 = 6'hf == cacheLine ? io_writeBlock[127:96] : cache_15_line_3; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1488 = 6'h10 == cacheLine ? io_writeBlock[127:96] : cache_16_line_3; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1489 = 6'h11 == cacheLine ? io_writeBlock[127:96] : cache_17_line_3; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1490 = 6'h12 == cacheLine ? io_writeBlock[127:96] : cache_18_line_3; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1491 = 6'h13 == cacheLine ? io_writeBlock[127:96] : cache_19_line_3; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1492 = 6'h14 == cacheLine ? io_writeBlock[127:96] : cache_20_line_3; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1493 = 6'h15 == cacheLine ? io_writeBlock[127:96] : cache_21_line_3; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1494 = 6'h16 == cacheLine ? io_writeBlock[127:96] : cache_22_line_3; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1495 = 6'h17 == cacheLine ? io_writeBlock[127:96] : cache_23_line_3; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1496 = 6'h18 == cacheLine ? io_writeBlock[127:96] : cache_24_line_3; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1497 = 6'h19 == cacheLine ? io_writeBlock[127:96] : cache_25_line_3; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1498 = 6'h1a == cacheLine ? io_writeBlock[127:96] : cache_26_line_3; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1499 = 6'h1b == cacheLine ? io_writeBlock[127:96] : cache_27_line_3; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1500 = 6'h1c == cacheLine ? io_writeBlock[127:96] : cache_28_line_3; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1501 = 6'h1d == cacheLine ? io_writeBlock[127:96] : cache_29_line_3; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1502 = 6'h1e == cacheLine ? io_writeBlock[127:96] : cache_30_line_3; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1503 = 6'h1f == cacheLine ? io_writeBlock[127:96] : cache_31_line_3; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1504 = 6'h20 == cacheLine ? io_writeBlock[127:96] : cache_32_line_3; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1505 = 6'h21 == cacheLine ? io_writeBlock[127:96] : cache_33_line_3; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1506 = 6'h22 == cacheLine ? io_writeBlock[127:96] : cache_34_line_3; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1507 = 6'h23 == cacheLine ? io_writeBlock[127:96] : cache_35_line_3; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1508 = 6'h24 == cacheLine ? io_writeBlock[127:96] : cache_36_line_3; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1509 = 6'h25 == cacheLine ? io_writeBlock[127:96] : cache_37_line_3; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1510 = 6'h26 == cacheLine ? io_writeBlock[127:96] : cache_38_line_3; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1511 = 6'h27 == cacheLine ? io_writeBlock[127:96] : cache_39_line_3; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1512 = 6'h28 == cacheLine ? io_writeBlock[127:96] : cache_40_line_3; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1513 = 6'h29 == cacheLine ? io_writeBlock[127:96] : cache_41_line_3; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1514 = 6'h2a == cacheLine ? io_writeBlock[127:96] : cache_42_line_3; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1515 = 6'h2b == cacheLine ? io_writeBlock[127:96] : cache_43_line_3; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1516 = 6'h2c == cacheLine ? io_writeBlock[127:96] : cache_44_line_3; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1517 = 6'h2d == cacheLine ? io_writeBlock[127:96] : cache_45_line_3; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1518 = 6'h2e == cacheLine ? io_writeBlock[127:96] : cache_46_line_3; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1519 = 6'h2f == cacheLine ? io_writeBlock[127:96] : cache_47_line_3; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1520 = 6'h30 == cacheLine ? io_writeBlock[127:96] : cache_48_line_3; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1521 = 6'h31 == cacheLine ? io_writeBlock[127:96] : cache_49_line_3; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1522 = 6'h32 == cacheLine ? io_writeBlock[127:96] : cache_50_line_3; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1523 = 6'h33 == cacheLine ? io_writeBlock[127:96] : cache_51_line_3; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1524 = 6'h34 == cacheLine ? io_writeBlock[127:96] : cache_52_line_3; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1525 = 6'h35 == cacheLine ? io_writeBlock[127:96] : cache_53_line_3; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1526 = 6'h36 == cacheLine ? io_writeBlock[127:96] : cache_54_line_3; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1527 = 6'h37 == cacheLine ? io_writeBlock[127:96] : cache_55_line_3; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1528 = 6'h38 == cacheLine ? io_writeBlock[127:96] : cache_56_line_3; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1529 = 6'h39 == cacheLine ? io_writeBlock[127:96] : cache_57_line_3; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1530 = 6'h3a == cacheLine ? io_writeBlock[127:96] : cache_58_line_3; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1531 = 6'h3b == cacheLine ? io_writeBlock[127:96] : cache_59_line_3; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1532 = 6'h3c == cacheLine ? io_writeBlock[127:96] : cache_60_line_3; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1533 = 6'h3d == cacheLine ? io_writeBlock[127:96] : cache_61_line_3; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1534 = 6'h3e == cacheLine ? io_writeBlock[127:96] : cache_62_line_3; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1535 = 6'h3f == cacheLine ? io_writeBlock[127:96] : cache_63_line_3; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1536 = 6'h0 == cacheLine ? io_writeBlock[159:128] : cache_0_line_4; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1537 = 6'h1 == cacheLine ? io_writeBlock[159:128] : cache_1_line_4; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1538 = 6'h2 == cacheLine ? io_writeBlock[159:128] : cache_2_line_4; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1539 = 6'h3 == cacheLine ? io_writeBlock[159:128] : cache_3_line_4; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1540 = 6'h4 == cacheLine ? io_writeBlock[159:128] : cache_4_line_4; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1541 = 6'h5 == cacheLine ? io_writeBlock[159:128] : cache_5_line_4; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1542 = 6'h6 == cacheLine ? io_writeBlock[159:128] : cache_6_line_4; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1543 = 6'h7 == cacheLine ? io_writeBlock[159:128] : cache_7_line_4; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1544 = 6'h8 == cacheLine ? io_writeBlock[159:128] : cache_8_line_4; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1545 = 6'h9 == cacheLine ? io_writeBlock[159:128] : cache_9_line_4; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1546 = 6'ha == cacheLine ? io_writeBlock[159:128] : cache_10_line_4; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1547 = 6'hb == cacheLine ? io_writeBlock[159:128] : cache_11_line_4; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1548 = 6'hc == cacheLine ? io_writeBlock[159:128] : cache_12_line_4; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1549 = 6'hd == cacheLine ? io_writeBlock[159:128] : cache_13_line_4; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1550 = 6'he == cacheLine ? io_writeBlock[159:128] : cache_14_line_4; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1551 = 6'hf == cacheLine ? io_writeBlock[159:128] : cache_15_line_4; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1552 = 6'h10 == cacheLine ? io_writeBlock[159:128] : cache_16_line_4; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1553 = 6'h11 == cacheLine ? io_writeBlock[159:128] : cache_17_line_4; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1554 = 6'h12 == cacheLine ? io_writeBlock[159:128] : cache_18_line_4; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1555 = 6'h13 == cacheLine ? io_writeBlock[159:128] : cache_19_line_4; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1556 = 6'h14 == cacheLine ? io_writeBlock[159:128] : cache_20_line_4; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1557 = 6'h15 == cacheLine ? io_writeBlock[159:128] : cache_21_line_4; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1558 = 6'h16 == cacheLine ? io_writeBlock[159:128] : cache_22_line_4; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1559 = 6'h17 == cacheLine ? io_writeBlock[159:128] : cache_23_line_4; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1560 = 6'h18 == cacheLine ? io_writeBlock[159:128] : cache_24_line_4; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1561 = 6'h19 == cacheLine ? io_writeBlock[159:128] : cache_25_line_4; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1562 = 6'h1a == cacheLine ? io_writeBlock[159:128] : cache_26_line_4; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1563 = 6'h1b == cacheLine ? io_writeBlock[159:128] : cache_27_line_4; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1564 = 6'h1c == cacheLine ? io_writeBlock[159:128] : cache_28_line_4; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1565 = 6'h1d == cacheLine ? io_writeBlock[159:128] : cache_29_line_4; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1566 = 6'h1e == cacheLine ? io_writeBlock[159:128] : cache_30_line_4; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1567 = 6'h1f == cacheLine ? io_writeBlock[159:128] : cache_31_line_4; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1568 = 6'h20 == cacheLine ? io_writeBlock[159:128] : cache_32_line_4; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1569 = 6'h21 == cacheLine ? io_writeBlock[159:128] : cache_33_line_4; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1570 = 6'h22 == cacheLine ? io_writeBlock[159:128] : cache_34_line_4; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1571 = 6'h23 == cacheLine ? io_writeBlock[159:128] : cache_35_line_4; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1572 = 6'h24 == cacheLine ? io_writeBlock[159:128] : cache_36_line_4; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1573 = 6'h25 == cacheLine ? io_writeBlock[159:128] : cache_37_line_4; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1574 = 6'h26 == cacheLine ? io_writeBlock[159:128] : cache_38_line_4; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1575 = 6'h27 == cacheLine ? io_writeBlock[159:128] : cache_39_line_4; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1576 = 6'h28 == cacheLine ? io_writeBlock[159:128] : cache_40_line_4; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1577 = 6'h29 == cacheLine ? io_writeBlock[159:128] : cache_41_line_4; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1578 = 6'h2a == cacheLine ? io_writeBlock[159:128] : cache_42_line_4; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1579 = 6'h2b == cacheLine ? io_writeBlock[159:128] : cache_43_line_4; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1580 = 6'h2c == cacheLine ? io_writeBlock[159:128] : cache_44_line_4; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1581 = 6'h2d == cacheLine ? io_writeBlock[159:128] : cache_45_line_4; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1582 = 6'h2e == cacheLine ? io_writeBlock[159:128] : cache_46_line_4; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1583 = 6'h2f == cacheLine ? io_writeBlock[159:128] : cache_47_line_4; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1584 = 6'h30 == cacheLine ? io_writeBlock[159:128] : cache_48_line_4; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1585 = 6'h31 == cacheLine ? io_writeBlock[159:128] : cache_49_line_4; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1586 = 6'h32 == cacheLine ? io_writeBlock[159:128] : cache_50_line_4; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1587 = 6'h33 == cacheLine ? io_writeBlock[159:128] : cache_51_line_4; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1588 = 6'h34 == cacheLine ? io_writeBlock[159:128] : cache_52_line_4; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1589 = 6'h35 == cacheLine ? io_writeBlock[159:128] : cache_53_line_4; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1590 = 6'h36 == cacheLine ? io_writeBlock[159:128] : cache_54_line_4; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1591 = 6'h37 == cacheLine ? io_writeBlock[159:128] : cache_55_line_4; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1592 = 6'h38 == cacheLine ? io_writeBlock[159:128] : cache_56_line_4; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1593 = 6'h39 == cacheLine ? io_writeBlock[159:128] : cache_57_line_4; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1594 = 6'h3a == cacheLine ? io_writeBlock[159:128] : cache_58_line_4; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1595 = 6'h3b == cacheLine ? io_writeBlock[159:128] : cache_59_line_4; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1596 = 6'h3c == cacheLine ? io_writeBlock[159:128] : cache_60_line_4; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1597 = 6'h3d == cacheLine ? io_writeBlock[159:128] : cache_61_line_4; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1598 = 6'h3e == cacheLine ? io_writeBlock[159:128] : cache_62_line_4; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1599 = 6'h3f == cacheLine ? io_writeBlock[159:128] : cache_63_line_4; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1600 = 6'h0 == cacheLine ? io_writeBlock[191:160] : cache_0_line_5; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1601 = 6'h1 == cacheLine ? io_writeBlock[191:160] : cache_1_line_5; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1602 = 6'h2 == cacheLine ? io_writeBlock[191:160] : cache_2_line_5; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1603 = 6'h3 == cacheLine ? io_writeBlock[191:160] : cache_3_line_5; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1604 = 6'h4 == cacheLine ? io_writeBlock[191:160] : cache_4_line_5; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1605 = 6'h5 == cacheLine ? io_writeBlock[191:160] : cache_5_line_5; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1606 = 6'h6 == cacheLine ? io_writeBlock[191:160] : cache_6_line_5; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1607 = 6'h7 == cacheLine ? io_writeBlock[191:160] : cache_7_line_5; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1608 = 6'h8 == cacheLine ? io_writeBlock[191:160] : cache_8_line_5; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1609 = 6'h9 == cacheLine ? io_writeBlock[191:160] : cache_9_line_5; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1610 = 6'ha == cacheLine ? io_writeBlock[191:160] : cache_10_line_5; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1611 = 6'hb == cacheLine ? io_writeBlock[191:160] : cache_11_line_5; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1612 = 6'hc == cacheLine ? io_writeBlock[191:160] : cache_12_line_5; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1613 = 6'hd == cacheLine ? io_writeBlock[191:160] : cache_13_line_5; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1614 = 6'he == cacheLine ? io_writeBlock[191:160] : cache_14_line_5; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1615 = 6'hf == cacheLine ? io_writeBlock[191:160] : cache_15_line_5; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1616 = 6'h10 == cacheLine ? io_writeBlock[191:160] : cache_16_line_5; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1617 = 6'h11 == cacheLine ? io_writeBlock[191:160] : cache_17_line_5; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1618 = 6'h12 == cacheLine ? io_writeBlock[191:160] : cache_18_line_5; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1619 = 6'h13 == cacheLine ? io_writeBlock[191:160] : cache_19_line_5; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1620 = 6'h14 == cacheLine ? io_writeBlock[191:160] : cache_20_line_5; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1621 = 6'h15 == cacheLine ? io_writeBlock[191:160] : cache_21_line_5; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1622 = 6'h16 == cacheLine ? io_writeBlock[191:160] : cache_22_line_5; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1623 = 6'h17 == cacheLine ? io_writeBlock[191:160] : cache_23_line_5; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1624 = 6'h18 == cacheLine ? io_writeBlock[191:160] : cache_24_line_5; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1625 = 6'h19 == cacheLine ? io_writeBlock[191:160] : cache_25_line_5; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1626 = 6'h1a == cacheLine ? io_writeBlock[191:160] : cache_26_line_5; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1627 = 6'h1b == cacheLine ? io_writeBlock[191:160] : cache_27_line_5; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1628 = 6'h1c == cacheLine ? io_writeBlock[191:160] : cache_28_line_5; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1629 = 6'h1d == cacheLine ? io_writeBlock[191:160] : cache_29_line_5; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1630 = 6'h1e == cacheLine ? io_writeBlock[191:160] : cache_30_line_5; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1631 = 6'h1f == cacheLine ? io_writeBlock[191:160] : cache_31_line_5; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1632 = 6'h20 == cacheLine ? io_writeBlock[191:160] : cache_32_line_5; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1633 = 6'h21 == cacheLine ? io_writeBlock[191:160] : cache_33_line_5; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1634 = 6'h22 == cacheLine ? io_writeBlock[191:160] : cache_34_line_5; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1635 = 6'h23 == cacheLine ? io_writeBlock[191:160] : cache_35_line_5; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1636 = 6'h24 == cacheLine ? io_writeBlock[191:160] : cache_36_line_5; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1637 = 6'h25 == cacheLine ? io_writeBlock[191:160] : cache_37_line_5; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1638 = 6'h26 == cacheLine ? io_writeBlock[191:160] : cache_38_line_5; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1639 = 6'h27 == cacheLine ? io_writeBlock[191:160] : cache_39_line_5; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1640 = 6'h28 == cacheLine ? io_writeBlock[191:160] : cache_40_line_5; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1641 = 6'h29 == cacheLine ? io_writeBlock[191:160] : cache_41_line_5; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1642 = 6'h2a == cacheLine ? io_writeBlock[191:160] : cache_42_line_5; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1643 = 6'h2b == cacheLine ? io_writeBlock[191:160] : cache_43_line_5; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1644 = 6'h2c == cacheLine ? io_writeBlock[191:160] : cache_44_line_5; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1645 = 6'h2d == cacheLine ? io_writeBlock[191:160] : cache_45_line_5; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1646 = 6'h2e == cacheLine ? io_writeBlock[191:160] : cache_46_line_5; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1647 = 6'h2f == cacheLine ? io_writeBlock[191:160] : cache_47_line_5; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1648 = 6'h30 == cacheLine ? io_writeBlock[191:160] : cache_48_line_5; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1649 = 6'h31 == cacheLine ? io_writeBlock[191:160] : cache_49_line_5; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1650 = 6'h32 == cacheLine ? io_writeBlock[191:160] : cache_50_line_5; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1651 = 6'h33 == cacheLine ? io_writeBlock[191:160] : cache_51_line_5; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1652 = 6'h34 == cacheLine ? io_writeBlock[191:160] : cache_52_line_5; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1653 = 6'h35 == cacheLine ? io_writeBlock[191:160] : cache_53_line_5; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1654 = 6'h36 == cacheLine ? io_writeBlock[191:160] : cache_54_line_5; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1655 = 6'h37 == cacheLine ? io_writeBlock[191:160] : cache_55_line_5; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1656 = 6'h38 == cacheLine ? io_writeBlock[191:160] : cache_56_line_5; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1657 = 6'h39 == cacheLine ? io_writeBlock[191:160] : cache_57_line_5; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1658 = 6'h3a == cacheLine ? io_writeBlock[191:160] : cache_58_line_5; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1659 = 6'h3b == cacheLine ? io_writeBlock[191:160] : cache_59_line_5; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1660 = 6'h3c == cacheLine ? io_writeBlock[191:160] : cache_60_line_5; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1661 = 6'h3d == cacheLine ? io_writeBlock[191:160] : cache_61_line_5; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1662 = 6'h3e == cacheLine ? io_writeBlock[191:160] : cache_62_line_5; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1663 = 6'h3f == cacheLine ? io_writeBlock[191:160] : cache_63_line_5; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1664 = 6'h0 == cacheLine ? io_writeBlock[223:192] : cache_0_line_6; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1665 = 6'h1 == cacheLine ? io_writeBlock[223:192] : cache_1_line_6; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1666 = 6'h2 == cacheLine ? io_writeBlock[223:192] : cache_2_line_6; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1667 = 6'h3 == cacheLine ? io_writeBlock[223:192] : cache_3_line_6; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1668 = 6'h4 == cacheLine ? io_writeBlock[223:192] : cache_4_line_6; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1669 = 6'h5 == cacheLine ? io_writeBlock[223:192] : cache_5_line_6; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1670 = 6'h6 == cacheLine ? io_writeBlock[223:192] : cache_6_line_6; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1671 = 6'h7 == cacheLine ? io_writeBlock[223:192] : cache_7_line_6; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1672 = 6'h8 == cacheLine ? io_writeBlock[223:192] : cache_8_line_6; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1673 = 6'h9 == cacheLine ? io_writeBlock[223:192] : cache_9_line_6; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1674 = 6'ha == cacheLine ? io_writeBlock[223:192] : cache_10_line_6; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1675 = 6'hb == cacheLine ? io_writeBlock[223:192] : cache_11_line_6; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1676 = 6'hc == cacheLine ? io_writeBlock[223:192] : cache_12_line_6; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1677 = 6'hd == cacheLine ? io_writeBlock[223:192] : cache_13_line_6; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1678 = 6'he == cacheLine ? io_writeBlock[223:192] : cache_14_line_6; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1679 = 6'hf == cacheLine ? io_writeBlock[223:192] : cache_15_line_6; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1680 = 6'h10 == cacheLine ? io_writeBlock[223:192] : cache_16_line_6; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1681 = 6'h11 == cacheLine ? io_writeBlock[223:192] : cache_17_line_6; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1682 = 6'h12 == cacheLine ? io_writeBlock[223:192] : cache_18_line_6; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1683 = 6'h13 == cacheLine ? io_writeBlock[223:192] : cache_19_line_6; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1684 = 6'h14 == cacheLine ? io_writeBlock[223:192] : cache_20_line_6; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1685 = 6'h15 == cacheLine ? io_writeBlock[223:192] : cache_21_line_6; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1686 = 6'h16 == cacheLine ? io_writeBlock[223:192] : cache_22_line_6; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1687 = 6'h17 == cacheLine ? io_writeBlock[223:192] : cache_23_line_6; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1688 = 6'h18 == cacheLine ? io_writeBlock[223:192] : cache_24_line_6; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1689 = 6'h19 == cacheLine ? io_writeBlock[223:192] : cache_25_line_6; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1690 = 6'h1a == cacheLine ? io_writeBlock[223:192] : cache_26_line_6; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1691 = 6'h1b == cacheLine ? io_writeBlock[223:192] : cache_27_line_6; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1692 = 6'h1c == cacheLine ? io_writeBlock[223:192] : cache_28_line_6; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1693 = 6'h1d == cacheLine ? io_writeBlock[223:192] : cache_29_line_6; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1694 = 6'h1e == cacheLine ? io_writeBlock[223:192] : cache_30_line_6; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1695 = 6'h1f == cacheLine ? io_writeBlock[223:192] : cache_31_line_6; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1696 = 6'h20 == cacheLine ? io_writeBlock[223:192] : cache_32_line_6; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1697 = 6'h21 == cacheLine ? io_writeBlock[223:192] : cache_33_line_6; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1698 = 6'h22 == cacheLine ? io_writeBlock[223:192] : cache_34_line_6; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1699 = 6'h23 == cacheLine ? io_writeBlock[223:192] : cache_35_line_6; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1700 = 6'h24 == cacheLine ? io_writeBlock[223:192] : cache_36_line_6; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1701 = 6'h25 == cacheLine ? io_writeBlock[223:192] : cache_37_line_6; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1702 = 6'h26 == cacheLine ? io_writeBlock[223:192] : cache_38_line_6; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1703 = 6'h27 == cacheLine ? io_writeBlock[223:192] : cache_39_line_6; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1704 = 6'h28 == cacheLine ? io_writeBlock[223:192] : cache_40_line_6; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1705 = 6'h29 == cacheLine ? io_writeBlock[223:192] : cache_41_line_6; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1706 = 6'h2a == cacheLine ? io_writeBlock[223:192] : cache_42_line_6; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1707 = 6'h2b == cacheLine ? io_writeBlock[223:192] : cache_43_line_6; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1708 = 6'h2c == cacheLine ? io_writeBlock[223:192] : cache_44_line_6; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1709 = 6'h2d == cacheLine ? io_writeBlock[223:192] : cache_45_line_6; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1710 = 6'h2e == cacheLine ? io_writeBlock[223:192] : cache_46_line_6; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1711 = 6'h2f == cacheLine ? io_writeBlock[223:192] : cache_47_line_6; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1712 = 6'h30 == cacheLine ? io_writeBlock[223:192] : cache_48_line_6; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1713 = 6'h31 == cacheLine ? io_writeBlock[223:192] : cache_49_line_6; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1714 = 6'h32 == cacheLine ? io_writeBlock[223:192] : cache_50_line_6; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1715 = 6'h33 == cacheLine ? io_writeBlock[223:192] : cache_51_line_6; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1716 = 6'h34 == cacheLine ? io_writeBlock[223:192] : cache_52_line_6; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1717 = 6'h35 == cacheLine ? io_writeBlock[223:192] : cache_53_line_6; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1718 = 6'h36 == cacheLine ? io_writeBlock[223:192] : cache_54_line_6; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1719 = 6'h37 == cacheLine ? io_writeBlock[223:192] : cache_55_line_6; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1720 = 6'h38 == cacheLine ? io_writeBlock[223:192] : cache_56_line_6; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1721 = 6'h39 == cacheLine ? io_writeBlock[223:192] : cache_57_line_6; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1722 = 6'h3a == cacheLine ? io_writeBlock[223:192] : cache_58_line_6; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1723 = 6'h3b == cacheLine ? io_writeBlock[223:192] : cache_59_line_6; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1724 = 6'h3c == cacheLine ? io_writeBlock[223:192] : cache_60_line_6; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1725 = 6'h3d == cacheLine ? io_writeBlock[223:192] : cache_61_line_6; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1726 = 6'h3e == cacheLine ? io_writeBlock[223:192] : cache_62_line_6; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1727 = 6'h3f == cacheLine ? io_writeBlock[223:192] : cache_63_line_6; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1728 = 6'h0 == cacheLine ? io_writeBlock[255:224] : cache_0_line_7; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1729 = 6'h1 == cacheLine ? io_writeBlock[255:224] : cache_1_line_7; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1730 = 6'h2 == cacheLine ? io_writeBlock[255:224] : cache_2_line_7; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1731 = 6'h3 == cacheLine ? io_writeBlock[255:224] : cache_3_line_7; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1732 = 6'h4 == cacheLine ? io_writeBlock[255:224] : cache_4_line_7; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1733 = 6'h5 == cacheLine ? io_writeBlock[255:224] : cache_5_line_7; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1734 = 6'h6 == cacheLine ? io_writeBlock[255:224] : cache_6_line_7; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1735 = 6'h7 == cacheLine ? io_writeBlock[255:224] : cache_7_line_7; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1736 = 6'h8 == cacheLine ? io_writeBlock[255:224] : cache_8_line_7; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1737 = 6'h9 == cacheLine ? io_writeBlock[255:224] : cache_9_line_7; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1738 = 6'ha == cacheLine ? io_writeBlock[255:224] : cache_10_line_7; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1739 = 6'hb == cacheLine ? io_writeBlock[255:224] : cache_11_line_7; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1740 = 6'hc == cacheLine ? io_writeBlock[255:224] : cache_12_line_7; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1741 = 6'hd == cacheLine ? io_writeBlock[255:224] : cache_13_line_7; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1742 = 6'he == cacheLine ? io_writeBlock[255:224] : cache_14_line_7; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1743 = 6'hf == cacheLine ? io_writeBlock[255:224] : cache_15_line_7; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1744 = 6'h10 == cacheLine ? io_writeBlock[255:224] : cache_16_line_7; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1745 = 6'h11 == cacheLine ? io_writeBlock[255:224] : cache_17_line_7; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1746 = 6'h12 == cacheLine ? io_writeBlock[255:224] : cache_18_line_7; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1747 = 6'h13 == cacheLine ? io_writeBlock[255:224] : cache_19_line_7; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1748 = 6'h14 == cacheLine ? io_writeBlock[255:224] : cache_20_line_7; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1749 = 6'h15 == cacheLine ? io_writeBlock[255:224] : cache_21_line_7; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1750 = 6'h16 == cacheLine ? io_writeBlock[255:224] : cache_22_line_7; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1751 = 6'h17 == cacheLine ? io_writeBlock[255:224] : cache_23_line_7; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1752 = 6'h18 == cacheLine ? io_writeBlock[255:224] : cache_24_line_7; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1753 = 6'h19 == cacheLine ? io_writeBlock[255:224] : cache_25_line_7; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1754 = 6'h1a == cacheLine ? io_writeBlock[255:224] : cache_26_line_7; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1755 = 6'h1b == cacheLine ? io_writeBlock[255:224] : cache_27_line_7; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1756 = 6'h1c == cacheLine ? io_writeBlock[255:224] : cache_28_line_7; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1757 = 6'h1d == cacheLine ? io_writeBlock[255:224] : cache_29_line_7; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1758 = 6'h1e == cacheLine ? io_writeBlock[255:224] : cache_30_line_7; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1759 = 6'h1f == cacheLine ? io_writeBlock[255:224] : cache_31_line_7; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1760 = 6'h20 == cacheLine ? io_writeBlock[255:224] : cache_32_line_7; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1761 = 6'h21 == cacheLine ? io_writeBlock[255:224] : cache_33_line_7; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1762 = 6'h22 == cacheLine ? io_writeBlock[255:224] : cache_34_line_7; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1763 = 6'h23 == cacheLine ? io_writeBlock[255:224] : cache_35_line_7; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1764 = 6'h24 == cacheLine ? io_writeBlock[255:224] : cache_36_line_7; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1765 = 6'h25 == cacheLine ? io_writeBlock[255:224] : cache_37_line_7; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1766 = 6'h26 == cacheLine ? io_writeBlock[255:224] : cache_38_line_7; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1767 = 6'h27 == cacheLine ? io_writeBlock[255:224] : cache_39_line_7; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1768 = 6'h28 == cacheLine ? io_writeBlock[255:224] : cache_40_line_7; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1769 = 6'h29 == cacheLine ? io_writeBlock[255:224] : cache_41_line_7; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1770 = 6'h2a == cacheLine ? io_writeBlock[255:224] : cache_42_line_7; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1771 = 6'h2b == cacheLine ? io_writeBlock[255:224] : cache_43_line_7; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1772 = 6'h2c == cacheLine ? io_writeBlock[255:224] : cache_44_line_7; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1773 = 6'h2d == cacheLine ? io_writeBlock[255:224] : cache_45_line_7; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1774 = 6'h2e == cacheLine ? io_writeBlock[255:224] : cache_46_line_7; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1775 = 6'h2f == cacheLine ? io_writeBlock[255:224] : cache_47_line_7; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1776 = 6'h30 == cacheLine ? io_writeBlock[255:224] : cache_48_line_7; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1777 = 6'h31 == cacheLine ? io_writeBlock[255:224] : cache_49_line_7; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1778 = 6'h32 == cacheLine ? io_writeBlock[255:224] : cache_50_line_7; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1779 = 6'h33 == cacheLine ? io_writeBlock[255:224] : cache_51_line_7; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1780 = 6'h34 == cacheLine ? io_writeBlock[255:224] : cache_52_line_7; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1781 = 6'h35 == cacheLine ? io_writeBlock[255:224] : cache_53_line_7; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1782 = 6'h36 == cacheLine ? io_writeBlock[255:224] : cache_54_line_7; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1783 = 6'h37 == cacheLine ? io_writeBlock[255:224] : cache_55_line_7; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1784 = 6'h38 == cacheLine ? io_writeBlock[255:224] : cache_56_line_7; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1785 = 6'h39 == cacheLine ? io_writeBlock[255:224] : cache_57_line_7; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1786 = 6'h3a == cacheLine ? io_writeBlock[255:224] : cache_58_line_7; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1787 = 6'h3b == cacheLine ? io_writeBlock[255:224] : cache_59_line_7; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1788 = 6'h3c == cacheLine ? io_writeBlock[255:224] : cache_60_line_7; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1789 = 6'h3d == cacheLine ? io_writeBlock[255:224] : cache_61_line_7; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1790 = 6'h3e == cacheLine ? io_writeBlock[255:224] : cache_62_line_7; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1791 = 6'h3f == cacheLine ? io_writeBlock[255:224] : cache_63_line_7; // @[Cache.scala 32:22 52:{34,34}]
  wire [31:0] _GEN_1920 = io_blockWriteEn ? _GEN_1280 : cache_0_line_0; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1921 = io_blockWriteEn ? _GEN_1281 : cache_1_line_0; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1922 = io_blockWriteEn ? _GEN_1282 : cache_2_line_0; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1923 = io_blockWriteEn ? _GEN_1283 : cache_3_line_0; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1924 = io_blockWriteEn ? _GEN_1284 : cache_4_line_0; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1925 = io_blockWriteEn ? _GEN_1285 : cache_5_line_0; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1926 = io_blockWriteEn ? _GEN_1286 : cache_6_line_0; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1927 = io_blockWriteEn ? _GEN_1287 : cache_7_line_0; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1928 = io_blockWriteEn ? _GEN_1288 : cache_8_line_0; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1929 = io_blockWriteEn ? _GEN_1289 : cache_9_line_0; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1930 = io_blockWriteEn ? _GEN_1290 : cache_10_line_0; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1931 = io_blockWriteEn ? _GEN_1291 : cache_11_line_0; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1932 = io_blockWriteEn ? _GEN_1292 : cache_12_line_0; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1933 = io_blockWriteEn ? _GEN_1293 : cache_13_line_0; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1934 = io_blockWriteEn ? _GEN_1294 : cache_14_line_0; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1935 = io_blockWriteEn ? _GEN_1295 : cache_15_line_0; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1936 = io_blockWriteEn ? _GEN_1296 : cache_16_line_0; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1937 = io_blockWriteEn ? _GEN_1297 : cache_17_line_0; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1938 = io_blockWriteEn ? _GEN_1298 : cache_18_line_0; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1939 = io_blockWriteEn ? _GEN_1299 : cache_19_line_0; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1940 = io_blockWriteEn ? _GEN_1300 : cache_20_line_0; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1941 = io_blockWriteEn ? _GEN_1301 : cache_21_line_0; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1942 = io_blockWriteEn ? _GEN_1302 : cache_22_line_0; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1943 = io_blockWriteEn ? _GEN_1303 : cache_23_line_0; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1944 = io_blockWriteEn ? _GEN_1304 : cache_24_line_0; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1945 = io_blockWriteEn ? _GEN_1305 : cache_25_line_0; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1946 = io_blockWriteEn ? _GEN_1306 : cache_26_line_0; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1947 = io_blockWriteEn ? _GEN_1307 : cache_27_line_0; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1948 = io_blockWriteEn ? _GEN_1308 : cache_28_line_0; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1949 = io_blockWriteEn ? _GEN_1309 : cache_29_line_0; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1950 = io_blockWriteEn ? _GEN_1310 : cache_30_line_0; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1951 = io_blockWriteEn ? _GEN_1311 : cache_31_line_0; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1952 = io_blockWriteEn ? _GEN_1312 : cache_32_line_0; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1953 = io_blockWriteEn ? _GEN_1313 : cache_33_line_0; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1954 = io_blockWriteEn ? _GEN_1314 : cache_34_line_0; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1955 = io_blockWriteEn ? _GEN_1315 : cache_35_line_0; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1956 = io_blockWriteEn ? _GEN_1316 : cache_36_line_0; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1957 = io_blockWriteEn ? _GEN_1317 : cache_37_line_0; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1958 = io_blockWriteEn ? _GEN_1318 : cache_38_line_0; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1959 = io_blockWriteEn ? _GEN_1319 : cache_39_line_0; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1960 = io_blockWriteEn ? _GEN_1320 : cache_40_line_0; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1961 = io_blockWriteEn ? _GEN_1321 : cache_41_line_0; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1962 = io_blockWriteEn ? _GEN_1322 : cache_42_line_0; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1963 = io_blockWriteEn ? _GEN_1323 : cache_43_line_0; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1964 = io_blockWriteEn ? _GEN_1324 : cache_44_line_0; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1965 = io_blockWriteEn ? _GEN_1325 : cache_45_line_0; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1966 = io_blockWriteEn ? _GEN_1326 : cache_46_line_0; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1967 = io_blockWriteEn ? _GEN_1327 : cache_47_line_0; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1968 = io_blockWriteEn ? _GEN_1328 : cache_48_line_0; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1969 = io_blockWriteEn ? _GEN_1329 : cache_49_line_0; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1970 = io_blockWriteEn ? _GEN_1330 : cache_50_line_0; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1971 = io_blockWriteEn ? _GEN_1331 : cache_51_line_0; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1972 = io_blockWriteEn ? _GEN_1332 : cache_52_line_0; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1973 = io_blockWriteEn ? _GEN_1333 : cache_53_line_0; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1974 = io_blockWriteEn ? _GEN_1334 : cache_54_line_0; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1975 = io_blockWriteEn ? _GEN_1335 : cache_55_line_0; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1976 = io_blockWriteEn ? _GEN_1336 : cache_56_line_0; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1977 = io_blockWriteEn ? _GEN_1337 : cache_57_line_0; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1978 = io_blockWriteEn ? _GEN_1338 : cache_58_line_0; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1979 = io_blockWriteEn ? _GEN_1339 : cache_59_line_0; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1980 = io_blockWriteEn ? _GEN_1340 : cache_60_line_0; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1981 = io_blockWriteEn ? _GEN_1341 : cache_61_line_0; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1982 = io_blockWriteEn ? _GEN_1342 : cache_62_line_0; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1983 = io_blockWriteEn ? _GEN_1343 : cache_63_line_0; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1984 = io_blockWriteEn ? _GEN_1344 : cache_0_line_1; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1985 = io_blockWriteEn ? _GEN_1345 : cache_1_line_1; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1986 = io_blockWriteEn ? _GEN_1346 : cache_2_line_1; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1987 = io_blockWriteEn ? _GEN_1347 : cache_3_line_1; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1988 = io_blockWriteEn ? _GEN_1348 : cache_4_line_1; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1989 = io_blockWriteEn ? _GEN_1349 : cache_5_line_1; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1990 = io_blockWriteEn ? _GEN_1350 : cache_6_line_1; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1991 = io_blockWriteEn ? _GEN_1351 : cache_7_line_1; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1992 = io_blockWriteEn ? _GEN_1352 : cache_8_line_1; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1993 = io_blockWriteEn ? _GEN_1353 : cache_9_line_1; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1994 = io_blockWriteEn ? _GEN_1354 : cache_10_line_1; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1995 = io_blockWriteEn ? _GEN_1355 : cache_11_line_1; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1996 = io_blockWriteEn ? _GEN_1356 : cache_12_line_1; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1997 = io_blockWriteEn ? _GEN_1357 : cache_13_line_1; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1998 = io_blockWriteEn ? _GEN_1358 : cache_14_line_1; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_1999 = io_blockWriteEn ? _GEN_1359 : cache_15_line_1; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2000 = io_blockWriteEn ? _GEN_1360 : cache_16_line_1; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2001 = io_blockWriteEn ? _GEN_1361 : cache_17_line_1; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2002 = io_blockWriteEn ? _GEN_1362 : cache_18_line_1; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2003 = io_blockWriteEn ? _GEN_1363 : cache_19_line_1; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2004 = io_blockWriteEn ? _GEN_1364 : cache_20_line_1; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2005 = io_blockWriteEn ? _GEN_1365 : cache_21_line_1; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2006 = io_blockWriteEn ? _GEN_1366 : cache_22_line_1; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2007 = io_blockWriteEn ? _GEN_1367 : cache_23_line_1; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2008 = io_blockWriteEn ? _GEN_1368 : cache_24_line_1; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2009 = io_blockWriteEn ? _GEN_1369 : cache_25_line_1; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2010 = io_blockWriteEn ? _GEN_1370 : cache_26_line_1; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2011 = io_blockWriteEn ? _GEN_1371 : cache_27_line_1; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2012 = io_blockWriteEn ? _GEN_1372 : cache_28_line_1; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2013 = io_blockWriteEn ? _GEN_1373 : cache_29_line_1; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2014 = io_blockWriteEn ? _GEN_1374 : cache_30_line_1; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2015 = io_blockWriteEn ? _GEN_1375 : cache_31_line_1; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2016 = io_blockWriteEn ? _GEN_1376 : cache_32_line_1; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2017 = io_blockWriteEn ? _GEN_1377 : cache_33_line_1; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2018 = io_blockWriteEn ? _GEN_1378 : cache_34_line_1; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2019 = io_blockWriteEn ? _GEN_1379 : cache_35_line_1; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2020 = io_blockWriteEn ? _GEN_1380 : cache_36_line_1; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2021 = io_blockWriteEn ? _GEN_1381 : cache_37_line_1; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2022 = io_blockWriteEn ? _GEN_1382 : cache_38_line_1; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2023 = io_blockWriteEn ? _GEN_1383 : cache_39_line_1; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2024 = io_blockWriteEn ? _GEN_1384 : cache_40_line_1; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2025 = io_blockWriteEn ? _GEN_1385 : cache_41_line_1; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2026 = io_blockWriteEn ? _GEN_1386 : cache_42_line_1; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2027 = io_blockWriteEn ? _GEN_1387 : cache_43_line_1; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2028 = io_blockWriteEn ? _GEN_1388 : cache_44_line_1; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2029 = io_blockWriteEn ? _GEN_1389 : cache_45_line_1; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2030 = io_blockWriteEn ? _GEN_1390 : cache_46_line_1; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2031 = io_blockWriteEn ? _GEN_1391 : cache_47_line_1; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2032 = io_blockWriteEn ? _GEN_1392 : cache_48_line_1; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2033 = io_blockWriteEn ? _GEN_1393 : cache_49_line_1; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2034 = io_blockWriteEn ? _GEN_1394 : cache_50_line_1; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2035 = io_blockWriteEn ? _GEN_1395 : cache_51_line_1; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2036 = io_blockWriteEn ? _GEN_1396 : cache_52_line_1; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2037 = io_blockWriteEn ? _GEN_1397 : cache_53_line_1; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2038 = io_blockWriteEn ? _GEN_1398 : cache_54_line_1; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2039 = io_blockWriteEn ? _GEN_1399 : cache_55_line_1; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2040 = io_blockWriteEn ? _GEN_1400 : cache_56_line_1; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2041 = io_blockWriteEn ? _GEN_1401 : cache_57_line_1; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2042 = io_blockWriteEn ? _GEN_1402 : cache_58_line_1; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2043 = io_blockWriteEn ? _GEN_1403 : cache_59_line_1; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2044 = io_blockWriteEn ? _GEN_1404 : cache_60_line_1; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2045 = io_blockWriteEn ? _GEN_1405 : cache_61_line_1; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2046 = io_blockWriteEn ? _GEN_1406 : cache_62_line_1; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2047 = io_blockWriteEn ? _GEN_1407 : cache_63_line_1; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2048 = io_blockWriteEn ? _GEN_1408 : cache_0_line_2; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2049 = io_blockWriteEn ? _GEN_1409 : cache_1_line_2; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2050 = io_blockWriteEn ? _GEN_1410 : cache_2_line_2; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2051 = io_blockWriteEn ? _GEN_1411 : cache_3_line_2; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2052 = io_blockWriteEn ? _GEN_1412 : cache_4_line_2; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2053 = io_blockWriteEn ? _GEN_1413 : cache_5_line_2; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2054 = io_blockWriteEn ? _GEN_1414 : cache_6_line_2; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2055 = io_blockWriteEn ? _GEN_1415 : cache_7_line_2; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2056 = io_blockWriteEn ? _GEN_1416 : cache_8_line_2; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2057 = io_blockWriteEn ? _GEN_1417 : cache_9_line_2; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2058 = io_blockWriteEn ? _GEN_1418 : cache_10_line_2; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2059 = io_blockWriteEn ? _GEN_1419 : cache_11_line_2; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2060 = io_blockWriteEn ? _GEN_1420 : cache_12_line_2; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2061 = io_blockWriteEn ? _GEN_1421 : cache_13_line_2; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2062 = io_blockWriteEn ? _GEN_1422 : cache_14_line_2; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2063 = io_blockWriteEn ? _GEN_1423 : cache_15_line_2; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2064 = io_blockWriteEn ? _GEN_1424 : cache_16_line_2; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2065 = io_blockWriteEn ? _GEN_1425 : cache_17_line_2; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2066 = io_blockWriteEn ? _GEN_1426 : cache_18_line_2; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2067 = io_blockWriteEn ? _GEN_1427 : cache_19_line_2; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2068 = io_blockWriteEn ? _GEN_1428 : cache_20_line_2; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2069 = io_blockWriteEn ? _GEN_1429 : cache_21_line_2; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2070 = io_blockWriteEn ? _GEN_1430 : cache_22_line_2; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2071 = io_blockWriteEn ? _GEN_1431 : cache_23_line_2; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2072 = io_blockWriteEn ? _GEN_1432 : cache_24_line_2; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2073 = io_blockWriteEn ? _GEN_1433 : cache_25_line_2; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2074 = io_blockWriteEn ? _GEN_1434 : cache_26_line_2; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2075 = io_blockWriteEn ? _GEN_1435 : cache_27_line_2; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2076 = io_blockWriteEn ? _GEN_1436 : cache_28_line_2; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2077 = io_blockWriteEn ? _GEN_1437 : cache_29_line_2; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2078 = io_blockWriteEn ? _GEN_1438 : cache_30_line_2; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2079 = io_blockWriteEn ? _GEN_1439 : cache_31_line_2; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2080 = io_blockWriteEn ? _GEN_1440 : cache_32_line_2; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2081 = io_blockWriteEn ? _GEN_1441 : cache_33_line_2; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2082 = io_blockWriteEn ? _GEN_1442 : cache_34_line_2; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2083 = io_blockWriteEn ? _GEN_1443 : cache_35_line_2; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2084 = io_blockWriteEn ? _GEN_1444 : cache_36_line_2; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2085 = io_blockWriteEn ? _GEN_1445 : cache_37_line_2; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2086 = io_blockWriteEn ? _GEN_1446 : cache_38_line_2; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2087 = io_blockWriteEn ? _GEN_1447 : cache_39_line_2; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2088 = io_blockWriteEn ? _GEN_1448 : cache_40_line_2; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2089 = io_blockWriteEn ? _GEN_1449 : cache_41_line_2; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2090 = io_blockWriteEn ? _GEN_1450 : cache_42_line_2; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2091 = io_blockWriteEn ? _GEN_1451 : cache_43_line_2; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2092 = io_blockWriteEn ? _GEN_1452 : cache_44_line_2; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2093 = io_blockWriteEn ? _GEN_1453 : cache_45_line_2; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2094 = io_blockWriteEn ? _GEN_1454 : cache_46_line_2; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2095 = io_blockWriteEn ? _GEN_1455 : cache_47_line_2; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2096 = io_blockWriteEn ? _GEN_1456 : cache_48_line_2; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2097 = io_blockWriteEn ? _GEN_1457 : cache_49_line_2; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2098 = io_blockWriteEn ? _GEN_1458 : cache_50_line_2; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2099 = io_blockWriteEn ? _GEN_1459 : cache_51_line_2; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2100 = io_blockWriteEn ? _GEN_1460 : cache_52_line_2; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2101 = io_blockWriteEn ? _GEN_1461 : cache_53_line_2; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2102 = io_blockWriteEn ? _GEN_1462 : cache_54_line_2; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2103 = io_blockWriteEn ? _GEN_1463 : cache_55_line_2; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2104 = io_blockWriteEn ? _GEN_1464 : cache_56_line_2; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2105 = io_blockWriteEn ? _GEN_1465 : cache_57_line_2; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2106 = io_blockWriteEn ? _GEN_1466 : cache_58_line_2; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2107 = io_blockWriteEn ? _GEN_1467 : cache_59_line_2; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2108 = io_blockWriteEn ? _GEN_1468 : cache_60_line_2; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2109 = io_blockWriteEn ? _GEN_1469 : cache_61_line_2; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2110 = io_blockWriteEn ? _GEN_1470 : cache_62_line_2; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2111 = io_blockWriteEn ? _GEN_1471 : cache_63_line_2; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2112 = io_blockWriteEn ? _GEN_1472 : cache_0_line_3; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2113 = io_blockWriteEn ? _GEN_1473 : cache_1_line_3; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2114 = io_blockWriteEn ? _GEN_1474 : cache_2_line_3; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2115 = io_blockWriteEn ? _GEN_1475 : cache_3_line_3; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2116 = io_blockWriteEn ? _GEN_1476 : cache_4_line_3; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2117 = io_blockWriteEn ? _GEN_1477 : cache_5_line_3; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2118 = io_blockWriteEn ? _GEN_1478 : cache_6_line_3; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2119 = io_blockWriteEn ? _GEN_1479 : cache_7_line_3; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2120 = io_blockWriteEn ? _GEN_1480 : cache_8_line_3; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2121 = io_blockWriteEn ? _GEN_1481 : cache_9_line_3; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2122 = io_blockWriteEn ? _GEN_1482 : cache_10_line_3; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2123 = io_blockWriteEn ? _GEN_1483 : cache_11_line_3; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2124 = io_blockWriteEn ? _GEN_1484 : cache_12_line_3; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2125 = io_blockWriteEn ? _GEN_1485 : cache_13_line_3; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2126 = io_blockWriteEn ? _GEN_1486 : cache_14_line_3; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2127 = io_blockWriteEn ? _GEN_1487 : cache_15_line_3; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2128 = io_blockWriteEn ? _GEN_1488 : cache_16_line_3; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2129 = io_blockWriteEn ? _GEN_1489 : cache_17_line_3; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2130 = io_blockWriteEn ? _GEN_1490 : cache_18_line_3; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2131 = io_blockWriteEn ? _GEN_1491 : cache_19_line_3; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2132 = io_blockWriteEn ? _GEN_1492 : cache_20_line_3; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2133 = io_blockWriteEn ? _GEN_1493 : cache_21_line_3; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2134 = io_blockWriteEn ? _GEN_1494 : cache_22_line_3; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2135 = io_blockWriteEn ? _GEN_1495 : cache_23_line_3; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2136 = io_blockWriteEn ? _GEN_1496 : cache_24_line_3; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2137 = io_blockWriteEn ? _GEN_1497 : cache_25_line_3; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2138 = io_blockWriteEn ? _GEN_1498 : cache_26_line_3; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2139 = io_blockWriteEn ? _GEN_1499 : cache_27_line_3; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2140 = io_blockWriteEn ? _GEN_1500 : cache_28_line_3; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2141 = io_blockWriteEn ? _GEN_1501 : cache_29_line_3; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2142 = io_blockWriteEn ? _GEN_1502 : cache_30_line_3; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2143 = io_blockWriteEn ? _GEN_1503 : cache_31_line_3; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2144 = io_blockWriteEn ? _GEN_1504 : cache_32_line_3; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2145 = io_blockWriteEn ? _GEN_1505 : cache_33_line_3; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2146 = io_blockWriteEn ? _GEN_1506 : cache_34_line_3; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2147 = io_blockWriteEn ? _GEN_1507 : cache_35_line_3; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2148 = io_blockWriteEn ? _GEN_1508 : cache_36_line_3; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2149 = io_blockWriteEn ? _GEN_1509 : cache_37_line_3; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2150 = io_blockWriteEn ? _GEN_1510 : cache_38_line_3; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2151 = io_blockWriteEn ? _GEN_1511 : cache_39_line_3; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2152 = io_blockWriteEn ? _GEN_1512 : cache_40_line_3; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2153 = io_blockWriteEn ? _GEN_1513 : cache_41_line_3; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2154 = io_blockWriteEn ? _GEN_1514 : cache_42_line_3; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2155 = io_blockWriteEn ? _GEN_1515 : cache_43_line_3; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2156 = io_blockWriteEn ? _GEN_1516 : cache_44_line_3; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2157 = io_blockWriteEn ? _GEN_1517 : cache_45_line_3; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2158 = io_blockWriteEn ? _GEN_1518 : cache_46_line_3; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2159 = io_blockWriteEn ? _GEN_1519 : cache_47_line_3; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2160 = io_blockWriteEn ? _GEN_1520 : cache_48_line_3; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2161 = io_blockWriteEn ? _GEN_1521 : cache_49_line_3; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2162 = io_blockWriteEn ? _GEN_1522 : cache_50_line_3; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2163 = io_blockWriteEn ? _GEN_1523 : cache_51_line_3; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2164 = io_blockWriteEn ? _GEN_1524 : cache_52_line_3; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2165 = io_blockWriteEn ? _GEN_1525 : cache_53_line_3; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2166 = io_blockWriteEn ? _GEN_1526 : cache_54_line_3; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2167 = io_blockWriteEn ? _GEN_1527 : cache_55_line_3; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2168 = io_blockWriteEn ? _GEN_1528 : cache_56_line_3; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2169 = io_blockWriteEn ? _GEN_1529 : cache_57_line_3; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2170 = io_blockWriteEn ? _GEN_1530 : cache_58_line_3; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2171 = io_blockWriteEn ? _GEN_1531 : cache_59_line_3; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2172 = io_blockWriteEn ? _GEN_1532 : cache_60_line_3; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2173 = io_blockWriteEn ? _GEN_1533 : cache_61_line_3; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2174 = io_blockWriteEn ? _GEN_1534 : cache_62_line_3; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2175 = io_blockWriteEn ? _GEN_1535 : cache_63_line_3; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2176 = io_blockWriteEn ? _GEN_1536 : cache_0_line_4; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2177 = io_blockWriteEn ? _GEN_1537 : cache_1_line_4; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2178 = io_blockWriteEn ? _GEN_1538 : cache_2_line_4; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2179 = io_blockWriteEn ? _GEN_1539 : cache_3_line_4; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2180 = io_blockWriteEn ? _GEN_1540 : cache_4_line_4; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2181 = io_blockWriteEn ? _GEN_1541 : cache_5_line_4; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2182 = io_blockWriteEn ? _GEN_1542 : cache_6_line_4; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2183 = io_blockWriteEn ? _GEN_1543 : cache_7_line_4; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2184 = io_blockWriteEn ? _GEN_1544 : cache_8_line_4; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2185 = io_blockWriteEn ? _GEN_1545 : cache_9_line_4; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2186 = io_blockWriteEn ? _GEN_1546 : cache_10_line_4; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2187 = io_blockWriteEn ? _GEN_1547 : cache_11_line_4; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2188 = io_blockWriteEn ? _GEN_1548 : cache_12_line_4; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2189 = io_blockWriteEn ? _GEN_1549 : cache_13_line_4; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2190 = io_blockWriteEn ? _GEN_1550 : cache_14_line_4; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2191 = io_blockWriteEn ? _GEN_1551 : cache_15_line_4; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2192 = io_blockWriteEn ? _GEN_1552 : cache_16_line_4; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2193 = io_blockWriteEn ? _GEN_1553 : cache_17_line_4; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2194 = io_blockWriteEn ? _GEN_1554 : cache_18_line_4; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2195 = io_blockWriteEn ? _GEN_1555 : cache_19_line_4; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2196 = io_blockWriteEn ? _GEN_1556 : cache_20_line_4; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2197 = io_blockWriteEn ? _GEN_1557 : cache_21_line_4; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2198 = io_blockWriteEn ? _GEN_1558 : cache_22_line_4; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2199 = io_blockWriteEn ? _GEN_1559 : cache_23_line_4; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2200 = io_blockWriteEn ? _GEN_1560 : cache_24_line_4; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2201 = io_blockWriteEn ? _GEN_1561 : cache_25_line_4; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2202 = io_blockWriteEn ? _GEN_1562 : cache_26_line_4; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2203 = io_blockWriteEn ? _GEN_1563 : cache_27_line_4; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2204 = io_blockWriteEn ? _GEN_1564 : cache_28_line_4; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2205 = io_blockWriteEn ? _GEN_1565 : cache_29_line_4; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2206 = io_blockWriteEn ? _GEN_1566 : cache_30_line_4; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2207 = io_blockWriteEn ? _GEN_1567 : cache_31_line_4; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2208 = io_blockWriteEn ? _GEN_1568 : cache_32_line_4; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2209 = io_blockWriteEn ? _GEN_1569 : cache_33_line_4; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2210 = io_blockWriteEn ? _GEN_1570 : cache_34_line_4; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2211 = io_blockWriteEn ? _GEN_1571 : cache_35_line_4; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2212 = io_blockWriteEn ? _GEN_1572 : cache_36_line_4; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2213 = io_blockWriteEn ? _GEN_1573 : cache_37_line_4; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2214 = io_blockWriteEn ? _GEN_1574 : cache_38_line_4; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2215 = io_blockWriteEn ? _GEN_1575 : cache_39_line_4; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2216 = io_blockWriteEn ? _GEN_1576 : cache_40_line_4; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2217 = io_blockWriteEn ? _GEN_1577 : cache_41_line_4; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2218 = io_blockWriteEn ? _GEN_1578 : cache_42_line_4; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2219 = io_blockWriteEn ? _GEN_1579 : cache_43_line_4; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2220 = io_blockWriteEn ? _GEN_1580 : cache_44_line_4; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2221 = io_blockWriteEn ? _GEN_1581 : cache_45_line_4; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2222 = io_blockWriteEn ? _GEN_1582 : cache_46_line_4; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2223 = io_blockWriteEn ? _GEN_1583 : cache_47_line_4; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2224 = io_blockWriteEn ? _GEN_1584 : cache_48_line_4; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2225 = io_blockWriteEn ? _GEN_1585 : cache_49_line_4; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2226 = io_blockWriteEn ? _GEN_1586 : cache_50_line_4; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2227 = io_blockWriteEn ? _GEN_1587 : cache_51_line_4; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2228 = io_blockWriteEn ? _GEN_1588 : cache_52_line_4; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2229 = io_blockWriteEn ? _GEN_1589 : cache_53_line_4; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2230 = io_blockWriteEn ? _GEN_1590 : cache_54_line_4; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2231 = io_blockWriteEn ? _GEN_1591 : cache_55_line_4; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2232 = io_blockWriteEn ? _GEN_1592 : cache_56_line_4; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2233 = io_blockWriteEn ? _GEN_1593 : cache_57_line_4; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2234 = io_blockWriteEn ? _GEN_1594 : cache_58_line_4; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2235 = io_blockWriteEn ? _GEN_1595 : cache_59_line_4; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2236 = io_blockWriteEn ? _GEN_1596 : cache_60_line_4; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2237 = io_blockWriteEn ? _GEN_1597 : cache_61_line_4; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2238 = io_blockWriteEn ? _GEN_1598 : cache_62_line_4; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2239 = io_blockWriteEn ? _GEN_1599 : cache_63_line_4; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2240 = io_blockWriteEn ? _GEN_1600 : cache_0_line_5; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2241 = io_blockWriteEn ? _GEN_1601 : cache_1_line_5; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2242 = io_blockWriteEn ? _GEN_1602 : cache_2_line_5; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2243 = io_blockWriteEn ? _GEN_1603 : cache_3_line_5; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2244 = io_blockWriteEn ? _GEN_1604 : cache_4_line_5; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2245 = io_blockWriteEn ? _GEN_1605 : cache_5_line_5; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2246 = io_blockWriteEn ? _GEN_1606 : cache_6_line_5; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2247 = io_blockWriteEn ? _GEN_1607 : cache_7_line_5; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2248 = io_blockWriteEn ? _GEN_1608 : cache_8_line_5; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2249 = io_blockWriteEn ? _GEN_1609 : cache_9_line_5; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2250 = io_blockWriteEn ? _GEN_1610 : cache_10_line_5; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2251 = io_blockWriteEn ? _GEN_1611 : cache_11_line_5; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2252 = io_blockWriteEn ? _GEN_1612 : cache_12_line_5; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2253 = io_blockWriteEn ? _GEN_1613 : cache_13_line_5; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2254 = io_blockWriteEn ? _GEN_1614 : cache_14_line_5; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2255 = io_blockWriteEn ? _GEN_1615 : cache_15_line_5; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2256 = io_blockWriteEn ? _GEN_1616 : cache_16_line_5; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2257 = io_blockWriteEn ? _GEN_1617 : cache_17_line_5; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2258 = io_blockWriteEn ? _GEN_1618 : cache_18_line_5; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2259 = io_blockWriteEn ? _GEN_1619 : cache_19_line_5; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2260 = io_blockWriteEn ? _GEN_1620 : cache_20_line_5; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2261 = io_blockWriteEn ? _GEN_1621 : cache_21_line_5; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2262 = io_blockWriteEn ? _GEN_1622 : cache_22_line_5; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2263 = io_blockWriteEn ? _GEN_1623 : cache_23_line_5; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2264 = io_blockWriteEn ? _GEN_1624 : cache_24_line_5; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2265 = io_blockWriteEn ? _GEN_1625 : cache_25_line_5; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2266 = io_blockWriteEn ? _GEN_1626 : cache_26_line_5; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2267 = io_blockWriteEn ? _GEN_1627 : cache_27_line_5; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2268 = io_blockWriteEn ? _GEN_1628 : cache_28_line_5; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2269 = io_blockWriteEn ? _GEN_1629 : cache_29_line_5; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2270 = io_blockWriteEn ? _GEN_1630 : cache_30_line_5; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2271 = io_blockWriteEn ? _GEN_1631 : cache_31_line_5; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2272 = io_blockWriteEn ? _GEN_1632 : cache_32_line_5; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2273 = io_blockWriteEn ? _GEN_1633 : cache_33_line_5; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2274 = io_blockWriteEn ? _GEN_1634 : cache_34_line_5; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2275 = io_blockWriteEn ? _GEN_1635 : cache_35_line_5; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2276 = io_blockWriteEn ? _GEN_1636 : cache_36_line_5; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2277 = io_blockWriteEn ? _GEN_1637 : cache_37_line_5; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2278 = io_blockWriteEn ? _GEN_1638 : cache_38_line_5; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2279 = io_blockWriteEn ? _GEN_1639 : cache_39_line_5; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2280 = io_blockWriteEn ? _GEN_1640 : cache_40_line_5; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2281 = io_blockWriteEn ? _GEN_1641 : cache_41_line_5; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2282 = io_blockWriteEn ? _GEN_1642 : cache_42_line_5; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2283 = io_blockWriteEn ? _GEN_1643 : cache_43_line_5; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2284 = io_blockWriteEn ? _GEN_1644 : cache_44_line_5; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2285 = io_blockWriteEn ? _GEN_1645 : cache_45_line_5; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2286 = io_blockWriteEn ? _GEN_1646 : cache_46_line_5; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2287 = io_blockWriteEn ? _GEN_1647 : cache_47_line_5; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2288 = io_blockWriteEn ? _GEN_1648 : cache_48_line_5; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2289 = io_blockWriteEn ? _GEN_1649 : cache_49_line_5; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2290 = io_blockWriteEn ? _GEN_1650 : cache_50_line_5; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2291 = io_blockWriteEn ? _GEN_1651 : cache_51_line_5; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2292 = io_blockWriteEn ? _GEN_1652 : cache_52_line_5; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2293 = io_blockWriteEn ? _GEN_1653 : cache_53_line_5; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2294 = io_blockWriteEn ? _GEN_1654 : cache_54_line_5; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2295 = io_blockWriteEn ? _GEN_1655 : cache_55_line_5; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2296 = io_blockWriteEn ? _GEN_1656 : cache_56_line_5; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2297 = io_blockWriteEn ? _GEN_1657 : cache_57_line_5; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2298 = io_blockWriteEn ? _GEN_1658 : cache_58_line_5; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2299 = io_blockWriteEn ? _GEN_1659 : cache_59_line_5; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2300 = io_blockWriteEn ? _GEN_1660 : cache_60_line_5; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2301 = io_blockWriteEn ? _GEN_1661 : cache_61_line_5; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2302 = io_blockWriteEn ? _GEN_1662 : cache_62_line_5; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2303 = io_blockWriteEn ? _GEN_1663 : cache_63_line_5; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2304 = io_blockWriteEn ? _GEN_1664 : cache_0_line_6; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2305 = io_blockWriteEn ? _GEN_1665 : cache_1_line_6; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2306 = io_blockWriteEn ? _GEN_1666 : cache_2_line_6; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2307 = io_blockWriteEn ? _GEN_1667 : cache_3_line_6; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2308 = io_blockWriteEn ? _GEN_1668 : cache_4_line_6; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2309 = io_blockWriteEn ? _GEN_1669 : cache_5_line_6; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2310 = io_blockWriteEn ? _GEN_1670 : cache_6_line_6; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2311 = io_blockWriteEn ? _GEN_1671 : cache_7_line_6; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2312 = io_blockWriteEn ? _GEN_1672 : cache_8_line_6; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2313 = io_blockWriteEn ? _GEN_1673 : cache_9_line_6; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2314 = io_blockWriteEn ? _GEN_1674 : cache_10_line_6; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2315 = io_blockWriteEn ? _GEN_1675 : cache_11_line_6; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2316 = io_blockWriteEn ? _GEN_1676 : cache_12_line_6; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2317 = io_blockWriteEn ? _GEN_1677 : cache_13_line_6; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2318 = io_blockWriteEn ? _GEN_1678 : cache_14_line_6; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2319 = io_blockWriteEn ? _GEN_1679 : cache_15_line_6; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2320 = io_blockWriteEn ? _GEN_1680 : cache_16_line_6; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2321 = io_blockWriteEn ? _GEN_1681 : cache_17_line_6; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2322 = io_blockWriteEn ? _GEN_1682 : cache_18_line_6; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2323 = io_blockWriteEn ? _GEN_1683 : cache_19_line_6; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2324 = io_blockWriteEn ? _GEN_1684 : cache_20_line_6; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2325 = io_blockWriteEn ? _GEN_1685 : cache_21_line_6; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2326 = io_blockWriteEn ? _GEN_1686 : cache_22_line_6; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2327 = io_blockWriteEn ? _GEN_1687 : cache_23_line_6; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2328 = io_blockWriteEn ? _GEN_1688 : cache_24_line_6; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2329 = io_blockWriteEn ? _GEN_1689 : cache_25_line_6; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2330 = io_blockWriteEn ? _GEN_1690 : cache_26_line_6; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2331 = io_blockWriteEn ? _GEN_1691 : cache_27_line_6; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2332 = io_blockWriteEn ? _GEN_1692 : cache_28_line_6; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2333 = io_blockWriteEn ? _GEN_1693 : cache_29_line_6; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2334 = io_blockWriteEn ? _GEN_1694 : cache_30_line_6; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2335 = io_blockWriteEn ? _GEN_1695 : cache_31_line_6; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2336 = io_blockWriteEn ? _GEN_1696 : cache_32_line_6; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2337 = io_blockWriteEn ? _GEN_1697 : cache_33_line_6; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2338 = io_blockWriteEn ? _GEN_1698 : cache_34_line_6; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2339 = io_blockWriteEn ? _GEN_1699 : cache_35_line_6; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2340 = io_blockWriteEn ? _GEN_1700 : cache_36_line_6; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2341 = io_blockWriteEn ? _GEN_1701 : cache_37_line_6; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2342 = io_blockWriteEn ? _GEN_1702 : cache_38_line_6; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2343 = io_blockWriteEn ? _GEN_1703 : cache_39_line_6; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2344 = io_blockWriteEn ? _GEN_1704 : cache_40_line_6; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2345 = io_blockWriteEn ? _GEN_1705 : cache_41_line_6; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2346 = io_blockWriteEn ? _GEN_1706 : cache_42_line_6; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2347 = io_blockWriteEn ? _GEN_1707 : cache_43_line_6; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2348 = io_blockWriteEn ? _GEN_1708 : cache_44_line_6; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2349 = io_blockWriteEn ? _GEN_1709 : cache_45_line_6; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2350 = io_blockWriteEn ? _GEN_1710 : cache_46_line_6; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2351 = io_blockWriteEn ? _GEN_1711 : cache_47_line_6; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2352 = io_blockWriteEn ? _GEN_1712 : cache_48_line_6; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2353 = io_blockWriteEn ? _GEN_1713 : cache_49_line_6; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2354 = io_blockWriteEn ? _GEN_1714 : cache_50_line_6; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2355 = io_blockWriteEn ? _GEN_1715 : cache_51_line_6; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2356 = io_blockWriteEn ? _GEN_1716 : cache_52_line_6; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2357 = io_blockWriteEn ? _GEN_1717 : cache_53_line_6; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2358 = io_blockWriteEn ? _GEN_1718 : cache_54_line_6; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2359 = io_blockWriteEn ? _GEN_1719 : cache_55_line_6; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2360 = io_blockWriteEn ? _GEN_1720 : cache_56_line_6; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2361 = io_blockWriteEn ? _GEN_1721 : cache_57_line_6; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2362 = io_blockWriteEn ? _GEN_1722 : cache_58_line_6; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2363 = io_blockWriteEn ? _GEN_1723 : cache_59_line_6; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2364 = io_blockWriteEn ? _GEN_1724 : cache_60_line_6; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2365 = io_blockWriteEn ? _GEN_1725 : cache_61_line_6; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2366 = io_blockWriteEn ? _GEN_1726 : cache_62_line_6; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2367 = io_blockWriteEn ? _GEN_1727 : cache_63_line_6; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2368 = io_blockWriteEn ? _GEN_1728 : cache_0_line_7; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2369 = io_blockWriteEn ? _GEN_1729 : cache_1_line_7; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2370 = io_blockWriteEn ? _GEN_1730 : cache_2_line_7; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2371 = io_blockWriteEn ? _GEN_1731 : cache_3_line_7; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2372 = io_blockWriteEn ? _GEN_1732 : cache_4_line_7; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2373 = io_blockWriteEn ? _GEN_1733 : cache_5_line_7; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2374 = io_blockWriteEn ? _GEN_1734 : cache_6_line_7; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2375 = io_blockWriteEn ? _GEN_1735 : cache_7_line_7; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2376 = io_blockWriteEn ? _GEN_1736 : cache_8_line_7; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2377 = io_blockWriteEn ? _GEN_1737 : cache_9_line_7; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2378 = io_blockWriteEn ? _GEN_1738 : cache_10_line_7; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2379 = io_blockWriteEn ? _GEN_1739 : cache_11_line_7; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2380 = io_blockWriteEn ? _GEN_1740 : cache_12_line_7; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2381 = io_blockWriteEn ? _GEN_1741 : cache_13_line_7; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2382 = io_blockWriteEn ? _GEN_1742 : cache_14_line_7; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2383 = io_blockWriteEn ? _GEN_1743 : cache_15_line_7; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2384 = io_blockWriteEn ? _GEN_1744 : cache_16_line_7; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2385 = io_blockWriteEn ? _GEN_1745 : cache_17_line_7; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2386 = io_blockWriteEn ? _GEN_1746 : cache_18_line_7; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2387 = io_blockWriteEn ? _GEN_1747 : cache_19_line_7; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2388 = io_blockWriteEn ? _GEN_1748 : cache_20_line_7; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2389 = io_blockWriteEn ? _GEN_1749 : cache_21_line_7; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2390 = io_blockWriteEn ? _GEN_1750 : cache_22_line_7; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2391 = io_blockWriteEn ? _GEN_1751 : cache_23_line_7; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2392 = io_blockWriteEn ? _GEN_1752 : cache_24_line_7; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2393 = io_blockWriteEn ? _GEN_1753 : cache_25_line_7; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2394 = io_blockWriteEn ? _GEN_1754 : cache_26_line_7; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2395 = io_blockWriteEn ? _GEN_1755 : cache_27_line_7; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2396 = io_blockWriteEn ? _GEN_1756 : cache_28_line_7; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2397 = io_blockWriteEn ? _GEN_1757 : cache_29_line_7; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2398 = io_blockWriteEn ? _GEN_1758 : cache_30_line_7; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2399 = io_blockWriteEn ? _GEN_1759 : cache_31_line_7; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2400 = io_blockWriteEn ? _GEN_1760 : cache_32_line_7; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2401 = io_blockWriteEn ? _GEN_1761 : cache_33_line_7; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2402 = io_blockWriteEn ? _GEN_1762 : cache_34_line_7; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2403 = io_blockWriteEn ? _GEN_1763 : cache_35_line_7; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2404 = io_blockWriteEn ? _GEN_1764 : cache_36_line_7; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2405 = io_blockWriteEn ? _GEN_1765 : cache_37_line_7; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2406 = io_blockWriteEn ? _GEN_1766 : cache_38_line_7; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2407 = io_blockWriteEn ? _GEN_1767 : cache_39_line_7; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2408 = io_blockWriteEn ? _GEN_1768 : cache_40_line_7; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2409 = io_blockWriteEn ? _GEN_1769 : cache_41_line_7; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2410 = io_blockWriteEn ? _GEN_1770 : cache_42_line_7; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2411 = io_blockWriteEn ? _GEN_1771 : cache_43_line_7; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2412 = io_blockWriteEn ? _GEN_1772 : cache_44_line_7; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2413 = io_blockWriteEn ? _GEN_1773 : cache_45_line_7; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2414 = io_blockWriteEn ? _GEN_1774 : cache_46_line_7; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2415 = io_blockWriteEn ? _GEN_1775 : cache_47_line_7; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2416 = io_blockWriteEn ? _GEN_1776 : cache_48_line_7; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2417 = io_blockWriteEn ? _GEN_1777 : cache_49_line_7; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2418 = io_blockWriteEn ? _GEN_1778 : cache_50_line_7; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2419 = io_blockWriteEn ? _GEN_1779 : cache_51_line_7; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2420 = io_blockWriteEn ? _GEN_1780 : cache_52_line_7; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2421 = io_blockWriteEn ? _GEN_1781 : cache_53_line_7; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2422 = io_blockWriteEn ? _GEN_1782 : cache_54_line_7; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2423 = io_blockWriteEn ? _GEN_1783 : cache_55_line_7; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2424 = io_blockWriteEn ? _GEN_1784 : cache_56_line_7; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2425 = io_blockWriteEn ? _GEN_1785 : cache_57_line_7; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2426 = io_blockWriteEn ? _GEN_1786 : cache_58_line_7; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2427 = io_blockWriteEn ? _GEN_1787 : cache_59_line_7; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2428 = io_blockWriteEn ? _GEN_1788 : cache_60_line_7; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2429 = io_blockWriteEn ? _GEN_1789 : cache_61_line_7; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2430 = io_blockWriteEn ? _GEN_1790 : cache_62_line_7; // @[Cache.scala 32:22 48:25]
  wire [31:0] _GEN_2431 = io_blockWriteEn ? _GEN_1791 : cache_63_line_7; // @[Cache.scala 32:22 48:25]
  wire [31:0] _cacheData_T_2 = {_GEN_639[31:8],io_cpuWriteData[7:0]}; // @[Cache.scala 62:34]
  wire [31:0] _cacheData_T_5 = {_GEN_639[31:16],io_cpuWriteData[15:0]}; // @[Cache.scala 65:35]
  wire [31:0] _GEN_2944 = 2'h2 == io_storeType ? io_cpuWriteData : 32'h0; // @[Cache.scala 60:26 68:19 57:30]
  wire [31:0] _GEN_2945 = 2'h1 == io_storeType ? _cacheData_T_5 : _GEN_2944; // @[Cache.scala 60:26 65:19]
  wire [31:0] _GEN_2946 = 2'h0 == io_storeType ? _cacheData_T_2 : _GEN_2945; // @[Cache.scala 60:26 62:19]
  assign io_cpuReadData = 6'h3f == cacheLine & 3'h7 == io_addrs[4:2] ? cache_63_line_7 : _GEN_638; // @[Cache.scala 40:{18,18}]
  assign io_bufferAddrs = addrsBuffer[10:0]; // @[Cache.scala 42:18]
  assign io_readBlock = dataBuffer; // @[Cache.scala 41:16]
  assign io_hit = _GEN_63 & tag == _GEN_127; // @[Cache.scala 39:32]
  always @(posedge clock) begin
    if (reset) begin // @[Cache.scala 32:22]
      cache_0_validBit <= 1'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      cache_0_validBit <= _GEN_1152;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_0_tag <= 5'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      if (6'h0 == cacheLine) begin // @[Cache.scala 50:26]
        cache_0_tag <= tag; // @[Cache.scala 50:26]
      end
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_0_line_0 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_3972 & _GEN_3987) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_0_line_0 <= _GEN_2946;
        end else begin
          cache_0_line_0 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_0_line_0 <= _GEN_1920;
      end
    end else begin
      cache_0_line_0 <= _GEN_1920;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_0_line_1 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_3972 & _GEN_3973) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_0_line_1 <= _GEN_2946;
        end else begin
          cache_0_line_1 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_0_line_1 <= _GEN_1984;
      end
    end else begin
      cache_0_line_1 <= _GEN_1984;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_0_line_2 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_3972 & _GEN_3975) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_0_line_2 <= _GEN_2946;
        end else begin
          cache_0_line_2 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_0_line_2 <= _GEN_2048;
      end
    end else begin
      cache_0_line_2 <= _GEN_2048;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_0_line_3 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_3972 & _GEN_3977) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_0_line_3 <= _GEN_2946;
        end else begin
          cache_0_line_3 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_0_line_3 <= _GEN_2112;
      end
    end else begin
      cache_0_line_3 <= _GEN_2112;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_0_line_4 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_3972 & _GEN_3979) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_0_line_4 <= _GEN_2946;
        end else begin
          cache_0_line_4 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_0_line_4 <= _GEN_2176;
      end
    end else begin
      cache_0_line_4 <= _GEN_2176;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_0_line_5 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_3972 & _GEN_3981) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_0_line_5 <= _GEN_2946;
        end else begin
          cache_0_line_5 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_0_line_5 <= _GEN_2240;
      end
    end else begin
      cache_0_line_5 <= _GEN_2240;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_0_line_6 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_3972 & _GEN_3983) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_0_line_6 <= _GEN_2946;
        end else begin
          cache_0_line_6 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_0_line_6 <= _GEN_2304;
      end
    end else begin
      cache_0_line_6 <= _GEN_2304;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_0_line_7 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_3972 & _GEN_3985) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_0_line_7 <= _GEN_2946;
        end else begin
          cache_0_line_7 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_0_line_7 <= _GEN_2368;
      end
    end else begin
      cache_0_line_7 <= _GEN_2368;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_1_validBit <= 1'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      cache_1_validBit <= _GEN_1153;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_1_tag <= 5'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      if (6'h1 == cacheLine) begin // @[Cache.scala 50:26]
        cache_1_tag <= tag; // @[Cache.scala 50:26]
      end
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_1_line_0 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_3986 & _GEN_3987) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_1_line_0 <= _GEN_2946;
        end else begin
          cache_1_line_0 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_1_line_0 <= _GEN_1921;
      end
    end else begin
      cache_1_line_0 <= _GEN_1921;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_1_line_1 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_3986 & _GEN_3973) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_1_line_1 <= _GEN_2946;
        end else begin
          cache_1_line_1 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_1_line_1 <= _GEN_1985;
      end
    end else begin
      cache_1_line_1 <= _GEN_1985;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_1_line_2 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_3986 & _GEN_3975) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_1_line_2 <= _GEN_2946;
        end else begin
          cache_1_line_2 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_1_line_2 <= _GEN_2049;
      end
    end else begin
      cache_1_line_2 <= _GEN_2049;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_1_line_3 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_3986 & _GEN_3977) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_1_line_3 <= _GEN_2946;
        end else begin
          cache_1_line_3 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_1_line_3 <= _GEN_2113;
      end
    end else begin
      cache_1_line_3 <= _GEN_2113;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_1_line_4 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_3986 & _GEN_3979) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_1_line_4 <= _GEN_2946;
        end else begin
          cache_1_line_4 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_1_line_4 <= _GEN_2177;
      end
    end else begin
      cache_1_line_4 <= _GEN_2177;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_1_line_5 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_3986 & _GEN_3981) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_1_line_5 <= _GEN_2946;
        end else begin
          cache_1_line_5 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_1_line_5 <= _GEN_2241;
      end
    end else begin
      cache_1_line_5 <= _GEN_2241;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_1_line_6 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_3986 & _GEN_3983) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_1_line_6 <= _GEN_2946;
        end else begin
          cache_1_line_6 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_1_line_6 <= _GEN_2305;
      end
    end else begin
      cache_1_line_6 <= _GEN_2305;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_1_line_7 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_3986 & _GEN_3985) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_1_line_7 <= _GEN_2946;
        end else begin
          cache_1_line_7 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_1_line_7 <= _GEN_2369;
      end
    end else begin
      cache_1_line_7 <= _GEN_2369;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_2_validBit <= 1'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      cache_2_validBit <= _GEN_1154;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_2_tag <= 5'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      if (6'h2 == cacheLine) begin // @[Cache.scala 50:26]
        cache_2_tag <= tag; // @[Cache.scala 50:26]
      end
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_2_line_0 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4002 & _GEN_3987) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_2_line_0 <= _GEN_2946;
        end else begin
          cache_2_line_0 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_2_line_0 <= _GEN_1922;
      end
    end else begin
      cache_2_line_0 <= _GEN_1922;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_2_line_1 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4002 & _GEN_3973) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_2_line_1 <= _GEN_2946;
        end else begin
          cache_2_line_1 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_2_line_1 <= _GEN_1986;
      end
    end else begin
      cache_2_line_1 <= _GEN_1986;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_2_line_2 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4002 & _GEN_3975) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_2_line_2 <= _GEN_2946;
        end else begin
          cache_2_line_2 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_2_line_2 <= _GEN_2050;
      end
    end else begin
      cache_2_line_2 <= _GEN_2050;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_2_line_3 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4002 & _GEN_3977) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_2_line_3 <= _GEN_2946;
        end else begin
          cache_2_line_3 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_2_line_3 <= _GEN_2114;
      end
    end else begin
      cache_2_line_3 <= _GEN_2114;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_2_line_4 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4002 & _GEN_3979) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_2_line_4 <= _GEN_2946;
        end else begin
          cache_2_line_4 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_2_line_4 <= _GEN_2178;
      end
    end else begin
      cache_2_line_4 <= _GEN_2178;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_2_line_5 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4002 & _GEN_3981) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_2_line_5 <= _GEN_2946;
        end else begin
          cache_2_line_5 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_2_line_5 <= _GEN_2242;
      end
    end else begin
      cache_2_line_5 <= _GEN_2242;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_2_line_6 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4002 & _GEN_3983) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_2_line_6 <= _GEN_2946;
        end else begin
          cache_2_line_6 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_2_line_6 <= _GEN_2306;
      end
    end else begin
      cache_2_line_6 <= _GEN_2306;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_2_line_7 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4002 & _GEN_3985) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_2_line_7 <= _GEN_2946;
        end else begin
          cache_2_line_7 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_2_line_7 <= _GEN_2370;
      end
    end else begin
      cache_2_line_7 <= _GEN_2370;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_3_validBit <= 1'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      cache_3_validBit <= _GEN_1155;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_3_tag <= 5'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      if (6'h3 == cacheLine) begin // @[Cache.scala 50:26]
        cache_3_tag <= tag; // @[Cache.scala 50:26]
      end
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_3_line_0 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4018 & _GEN_3987) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_3_line_0 <= _GEN_2946;
        end else begin
          cache_3_line_0 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_3_line_0 <= _GEN_1923;
      end
    end else begin
      cache_3_line_0 <= _GEN_1923;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_3_line_1 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4018 & _GEN_3973) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_3_line_1 <= _GEN_2946;
        end else begin
          cache_3_line_1 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_3_line_1 <= _GEN_1987;
      end
    end else begin
      cache_3_line_1 <= _GEN_1987;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_3_line_2 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4018 & _GEN_3975) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_3_line_2 <= _GEN_2946;
        end else begin
          cache_3_line_2 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_3_line_2 <= _GEN_2051;
      end
    end else begin
      cache_3_line_2 <= _GEN_2051;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_3_line_3 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4018 & _GEN_3977) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_3_line_3 <= _GEN_2946;
        end else begin
          cache_3_line_3 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_3_line_3 <= _GEN_2115;
      end
    end else begin
      cache_3_line_3 <= _GEN_2115;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_3_line_4 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4018 & _GEN_3979) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_3_line_4 <= _GEN_2946;
        end else begin
          cache_3_line_4 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_3_line_4 <= _GEN_2179;
      end
    end else begin
      cache_3_line_4 <= _GEN_2179;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_3_line_5 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4018 & _GEN_3981) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_3_line_5 <= _GEN_2946;
        end else begin
          cache_3_line_5 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_3_line_5 <= _GEN_2243;
      end
    end else begin
      cache_3_line_5 <= _GEN_2243;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_3_line_6 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4018 & _GEN_3983) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_3_line_6 <= _GEN_2946;
        end else begin
          cache_3_line_6 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_3_line_6 <= _GEN_2307;
      end
    end else begin
      cache_3_line_6 <= _GEN_2307;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_3_line_7 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4018 & _GEN_3985) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_3_line_7 <= _GEN_2946;
        end else begin
          cache_3_line_7 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_3_line_7 <= _GEN_2371;
      end
    end else begin
      cache_3_line_7 <= _GEN_2371;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_4_validBit <= 1'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      cache_4_validBit <= _GEN_1156;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_4_tag <= 5'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      if (6'h4 == cacheLine) begin // @[Cache.scala 50:26]
        cache_4_tag <= tag; // @[Cache.scala 50:26]
      end
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_4_line_0 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4034 & _GEN_3987) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_4_line_0 <= _GEN_2946;
        end else begin
          cache_4_line_0 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_4_line_0 <= _GEN_1924;
      end
    end else begin
      cache_4_line_0 <= _GEN_1924;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_4_line_1 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4034 & _GEN_3973) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_4_line_1 <= _GEN_2946;
        end else begin
          cache_4_line_1 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_4_line_1 <= _GEN_1988;
      end
    end else begin
      cache_4_line_1 <= _GEN_1988;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_4_line_2 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4034 & _GEN_3975) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_4_line_2 <= _GEN_2946;
        end else begin
          cache_4_line_2 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_4_line_2 <= _GEN_2052;
      end
    end else begin
      cache_4_line_2 <= _GEN_2052;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_4_line_3 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4034 & _GEN_3977) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_4_line_3 <= _GEN_2946;
        end else begin
          cache_4_line_3 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_4_line_3 <= _GEN_2116;
      end
    end else begin
      cache_4_line_3 <= _GEN_2116;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_4_line_4 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4034 & _GEN_3979) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_4_line_4 <= _GEN_2946;
        end else begin
          cache_4_line_4 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_4_line_4 <= _GEN_2180;
      end
    end else begin
      cache_4_line_4 <= _GEN_2180;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_4_line_5 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4034 & _GEN_3981) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_4_line_5 <= _GEN_2946;
        end else begin
          cache_4_line_5 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_4_line_5 <= _GEN_2244;
      end
    end else begin
      cache_4_line_5 <= _GEN_2244;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_4_line_6 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4034 & _GEN_3983) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_4_line_6 <= _GEN_2946;
        end else begin
          cache_4_line_6 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_4_line_6 <= _GEN_2308;
      end
    end else begin
      cache_4_line_6 <= _GEN_2308;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_4_line_7 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4034 & _GEN_3985) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_4_line_7 <= _GEN_2946;
        end else begin
          cache_4_line_7 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_4_line_7 <= _GEN_2372;
      end
    end else begin
      cache_4_line_7 <= _GEN_2372;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_5_validBit <= 1'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      cache_5_validBit <= _GEN_1157;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_5_tag <= 5'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      if (6'h5 == cacheLine) begin // @[Cache.scala 50:26]
        cache_5_tag <= tag; // @[Cache.scala 50:26]
      end
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_5_line_0 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4050 & _GEN_3987) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_5_line_0 <= _GEN_2946;
        end else begin
          cache_5_line_0 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_5_line_0 <= _GEN_1925;
      end
    end else begin
      cache_5_line_0 <= _GEN_1925;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_5_line_1 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4050 & _GEN_3973) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_5_line_1 <= _GEN_2946;
        end else begin
          cache_5_line_1 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_5_line_1 <= _GEN_1989;
      end
    end else begin
      cache_5_line_1 <= _GEN_1989;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_5_line_2 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4050 & _GEN_3975) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_5_line_2 <= _GEN_2946;
        end else begin
          cache_5_line_2 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_5_line_2 <= _GEN_2053;
      end
    end else begin
      cache_5_line_2 <= _GEN_2053;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_5_line_3 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4050 & _GEN_3977) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_5_line_3 <= _GEN_2946;
        end else begin
          cache_5_line_3 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_5_line_3 <= _GEN_2117;
      end
    end else begin
      cache_5_line_3 <= _GEN_2117;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_5_line_4 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4050 & _GEN_3979) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_5_line_4 <= _GEN_2946;
        end else begin
          cache_5_line_4 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_5_line_4 <= _GEN_2181;
      end
    end else begin
      cache_5_line_4 <= _GEN_2181;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_5_line_5 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4050 & _GEN_3981) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_5_line_5 <= _GEN_2946;
        end else begin
          cache_5_line_5 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_5_line_5 <= _GEN_2245;
      end
    end else begin
      cache_5_line_5 <= _GEN_2245;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_5_line_6 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4050 & _GEN_3983) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_5_line_6 <= _GEN_2946;
        end else begin
          cache_5_line_6 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_5_line_6 <= _GEN_2309;
      end
    end else begin
      cache_5_line_6 <= _GEN_2309;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_5_line_7 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4050 & _GEN_3985) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_5_line_7 <= _GEN_2946;
        end else begin
          cache_5_line_7 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_5_line_7 <= _GEN_2373;
      end
    end else begin
      cache_5_line_7 <= _GEN_2373;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_6_validBit <= 1'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      cache_6_validBit <= _GEN_1158;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_6_tag <= 5'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      if (6'h6 == cacheLine) begin // @[Cache.scala 50:26]
        cache_6_tag <= tag; // @[Cache.scala 50:26]
      end
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_6_line_0 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4066 & _GEN_3987) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_6_line_0 <= _GEN_2946;
        end else begin
          cache_6_line_0 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_6_line_0 <= _GEN_1926;
      end
    end else begin
      cache_6_line_0 <= _GEN_1926;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_6_line_1 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4066 & _GEN_3973) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_6_line_1 <= _GEN_2946;
        end else begin
          cache_6_line_1 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_6_line_1 <= _GEN_1990;
      end
    end else begin
      cache_6_line_1 <= _GEN_1990;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_6_line_2 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4066 & _GEN_3975) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_6_line_2 <= _GEN_2946;
        end else begin
          cache_6_line_2 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_6_line_2 <= _GEN_2054;
      end
    end else begin
      cache_6_line_2 <= _GEN_2054;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_6_line_3 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4066 & _GEN_3977) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_6_line_3 <= _GEN_2946;
        end else begin
          cache_6_line_3 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_6_line_3 <= _GEN_2118;
      end
    end else begin
      cache_6_line_3 <= _GEN_2118;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_6_line_4 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4066 & _GEN_3979) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_6_line_4 <= _GEN_2946;
        end else begin
          cache_6_line_4 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_6_line_4 <= _GEN_2182;
      end
    end else begin
      cache_6_line_4 <= _GEN_2182;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_6_line_5 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4066 & _GEN_3981) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_6_line_5 <= _GEN_2946;
        end else begin
          cache_6_line_5 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_6_line_5 <= _GEN_2246;
      end
    end else begin
      cache_6_line_5 <= _GEN_2246;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_6_line_6 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4066 & _GEN_3983) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_6_line_6 <= _GEN_2946;
        end else begin
          cache_6_line_6 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_6_line_6 <= _GEN_2310;
      end
    end else begin
      cache_6_line_6 <= _GEN_2310;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_6_line_7 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4066 & _GEN_3985) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_6_line_7 <= _GEN_2946;
        end else begin
          cache_6_line_7 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_6_line_7 <= _GEN_2374;
      end
    end else begin
      cache_6_line_7 <= _GEN_2374;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_7_validBit <= 1'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      cache_7_validBit <= _GEN_1159;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_7_tag <= 5'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      if (6'h7 == cacheLine) begin // @[Cache.scala 50:26]
        cache_7_tag <= tag; // @[Cache.scala 50:26]
      end
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_7_line_0 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4082 & _GEN_3987) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_7_line_0 <= _GEN_2946;
        end else begin
          cache_7_line_0 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_7_line_0 <= _GEN_1927;
      end
    end else begin
      cache_7_line_0 <= _GEN_1927;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_7_line_1 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4082 & _GEN_3973) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_7_line_1 <= _GEN_2946;
        end else begin
          cache_7_line_1 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_7_line_1 <= _GEN_1991;
      end
    end else begin
      cache_7_line_1 <= _GEN_1991;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_7_line_2 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4082 & _GEN_3975) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_7_line_2 <= _GEN_2946;
        end else begin
          cache_7_line_2 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_7_line_2 <= _GEN_2055;
      end
    end else begin
      cache_7_line_2 <= _GEN_2055;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_7_line_3 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4082 & _GEN_3977) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_7_line_3 <= _GEN_2946;
        end else begin
          cache_7_line_3 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_7_line_3 <= _GEN_2119;
      end
    end else begin
      cache_7_line_3 <= _GEN_2119;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_7_line_4 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4082 & _GEN_3979) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_7_line_4 <= _GEN_2946;
        end else begin
          cache_7_line_4 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_7_line_4 <= _GEN_2183;
      end
    end else begin
      cache_7_line_4 <= _GEN_2183;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_7_line_5 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4082 & _GEN_3981) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_7_line_5 <= _GEN_2946;
        end else begin
          cache_7_line_5 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_7_line_5 <= _GEN_2247;
      end
    end else begin
      cache_7_line_5 <= _GEN_2247;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_7_line_6 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4082 & _GEN_3983) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_7_line_6 <= _GEN_2946;
        end else begin
          cache_7_line_6 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_7_line_6 <= _GEN_2311;
      end
    end else begin
      cache_7_line_6 <= _GEN_2311;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_7_line_7 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4082 & _GEN_3985) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_7_line_7 <= _GEN_2946;
        end else begin
          cache_7_line_7 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_7_line_7 <= _GEN_2375;
      end
    end else begin
      cache_7_line_7 <= _GEN_2375;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_8_validBit <= 1'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      cache_8_validBit <= _GEN_1160;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_8_tag <= 5'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      if (6'h8 == cacheLine) begin // @[Cache.scala 50:26]
        cache_8_tag <= tag; // @[Cache.scala 50:26]
      end
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_8_line_0 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4098 & _GEN_3987) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_8_line_0 <= _GEN_2946;
        end else begin
          cache_8_line_0 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_8_line_0 <= _GEN_1928;
      end
    end else begin
      cache_8_line_0 <= _GEN_1928;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_8_line_1 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4098 & _GEN_3973) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_8_line_1 <= _GEN_2946;
        end else begin
          cache_8_line_1 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_8_line_1 <= _GEN_1992;
      end
    end else begin
      cache_8_line_1 <= _GEN_1992;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_8_line_2 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4098 & _GEN_3975) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_8_line_2 <= _GEN_2946;
        end else begin
          cache_8_line_2 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_8_line_2 <= _GEN_2056;
      end
    end else begin
      cache_8_line_2 <= _GEN_2056;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_8_line_3 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4098 & _GEN_3977) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_8_line_3 <= _GEN_2946;
        end else begin
          cache_8_line_3 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_8_line_3 <= _GEN_2120;
      end
    end else begin
      cache_8_line_3 <= _GEN_2120;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_8_line_4 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4098 & _GEN_3979) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_8_line_4 <= _GEN_2946;
        end else begin
          cache_8_line_4 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_8_line_4 <= _GEN_2184;
      end
    end else begin
      cache_8_line_4 <= _GEN_2184;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_8_line_5 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4098 & _GEN_3981) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_8_line_5 <= _GEN_2946;
        end else begin
          cache_8_line_5 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_8_line_5 <= _GEN_2248;
      end
    end else begin
      cache_8_line_5 <= _GEN_2248;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_8_line_6 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4098 & _GEN_3983) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_8_line_6 <= _GEN_2946;
        end else begin
          cache_8_line_6 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_8_line_6 <= _GEN_2312;
      end
    end else begin
      cache_8_line_6 <= _GEN_2312;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_8_line_7 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4098 & _GEN_3985) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_8_line_7 <= _GEN_2946;
        end else begin
          cache_8_line_7 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_8_line_7 <= _GEN_2376;
      end
    end else begin
      cache_8_line_7 <= _GEN_2376;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_9_validBit <= 1'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      cache_9_validBit <= _GEN_1161;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_9_tag <= 5'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      if (6'h9 == cacheLine) begin // @[Cache.scala 50:26]
        cache_9_tag <= tag; // @[Cache.scala 50:26]
      end
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_9_line_0 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4114 & _GEN_3987) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_9_line_0 <= _GEN_2946;
        end else begin
          cache_9_line_0 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_9_line_0 <= _GEN_1929;
      end
    end else begin
      cache_9_line_0 <= _GEN_1929;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_9_line_1 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4114 & _GEN_3973) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_9_line_1 <= _GEN_2946;
        end else begin
          cache_9_line_1 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_9_line_1 <= _GEN_1993;
      end
    end else begin
      cache_9_line_1 <= _GEN_1993;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_9_line_2 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4114 & _GEN_3975) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_9_line_2 <= _GEN_2946;
        end else begin
          cache_9_line_2 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_9_line_2 <= _GEN_2057;
      end
    end else begin
      cache_9_line_2 <= _GEN_2057;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_9_line_3 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4114 & _GEN_3977) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_9_line_3 <= _GEN_2946;
        end else begin
          cache_9_line_3 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_9_line_3 <= _GEN_2121;
      end
    end else begin
      cache_9_line_3 <= _GEN_2121;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_9_line_4 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4114 & _GEN_3979) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_9_line_4 <= _GEN_2946;
        end else begin
          cache_9_line_4 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_9_line_4 <= _GEN_2185;
      end
    end else begin
      cache_9_line_4 <= _GEN_2185;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_9_line_5 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4114 & _GEN_3981) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_9_line_5 <= _GEN_2946;
        end else begin
          cache_9_line_5 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_9_line_5 <= _GEN_2249;
      end
    end else begin
      cache_9_line_5 <= _GEN_2249;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_9_line_6 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4114 & _GEN_3983) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_9_line_6 <= _GEN_2946;
        end else begin
          cache_9_line_6 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_9_line_6 <= _GEN_2313;
      end
    end else begin
      cache_9_line_6 <= _GEN_2313;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_9_line_7 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4114 & _GEN_3985) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_9_line_7 <= _GEN_2946;
        end else begin
          cache_9_line_7 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_9_line_7 <= _GEN_2377;
      end
    end else begin
      cache_9_line_7 <= _GEN_2377;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_10_validBit <= 1'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      cache_10_validBit <= _GEN_1162;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_10_tag <= 5'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      if (6'ha == cacheLine) begin // @[Cache.scala 50:26]
        cache_10_tag <= tag; // @[Cache.scala 50:26]
      end
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_10_line_0 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4130 & _GEN_3987) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_10_line_0 <= _GEN_2946;
        end else begin
          cache_10_line_0 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_10_line_0 <= _GEN_1930;
      end
    end else begin
      cache_10_line_0 <= _GEN_1930;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_10_line_1 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4130 & _GEN_3973) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_10_line_1 <= _GEN_2946;
        end else begin
          cache_10_line_1 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_10_line_1 <= _GEN_1994;
      end
    end else begin
      cache_10_line_1 <= _GEN_1994;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_10_line_2 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4130 & _GEN_3975) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_10_line_2 <= _GEN_2946;
        end else begin
          cache_10_line_2 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_10_line_2 <= _GEN_2058;
      end
    end else begin
      cache_10_line_2 <= _GEN_2058;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_10_line_3 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4130 & _GEN_3977) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_10_line_3 <= _GEN_2946;
        end else begin
          cache_10_line_3 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_10_line_3 <= _GEN_2122;
      end
    end else begin
      cache_10_line_3 <= _GEN_2122;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_10_line_4 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4130 & _GEN_3979) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_10_line_4 <= _GEN_2946;
        end else begin
          cache_10_line_4 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_10_line_4 <= _GEN_2186;
      end
    end else begin
      cache_10_line_4 <= _GEN_2186;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_10_line_5 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4130 & _GEN_3981) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_10_line_5 <= _GEN_2946;
        end else begin
          cache_10_line_5 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_10_line_5 <= _GEN_2250;
      end
    end else begin
      cache_10_line_5 <= _GEN_2250;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_10_line_6 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4130 & _GEN_3983) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_10_line_6 <= _GEN_2946;
        end else begin
          cache_10_line_6 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_10_line_6 <= _GEN_2314;
      end
    end else begin
      cache_10_line_6 <= _GEN_2314;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_10_line_7 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4130 & _GEN_3985) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_10_line_7 <= _GEN_2946;
        end else begin
          cache_10_line_7 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_10_line_7 <= _GEN_2378;
      end
    end else begin
      cache_10_line_7 <= _GEN_2378;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_11_validBit <= 1'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      cache_11_validBit <= _GEN_1163;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_11_tag <= 5'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      if (6'hb == cacheLine) begin // @[Cache.scala 50:26]
        cache_11_tag <= tag; // @[Cache.scala 50:26]
      end
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_11_line_0 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4146 & _GEN_3987) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_11_line_0 <= _GEN_2946;
        end else begin
          cache_11_line_0 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_11_line_0 <= _GEN_1931;
      end
    end else begin
      cache_11_line_0 <= _GEN_1931;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_11_line_1 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4146 & _GEN_3973) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_11_line_1 <= _GEN_2946;
        end else begin
          cache_11_line_1 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_11_line_1 <= _GEN_1995;
      end
    end else begin
      cache_11_line_1 <= _GEN_1995;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_11_line_2 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4146 & _GEN_3975) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_11_line_2 <= _GEN_2946;
        end else begin
          cache_11_line_2 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_11_line_2 <= _GEN_2059;
      end
    end else begin
      cache_11_line_2 <= _GEN_2059;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_11_line_3 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4146 & _GEN_3977) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_11_line_3 <= _GEN_2946;
        end else begin
          cache_11_line_3 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_11_line_3 <= _GEN_2123;
      end
    end else begin
      cache_11_line_3 <= _GEN_2123;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_11_line_4 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4146 & _GEN_3979) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_11_line_4 <= _GEN_2946;
        end else begin
          cache_11_line_4 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_11_line_4 <= _GEN_2187;
      end
    end else begin
      cache_11_line_4 <= _GEN_2187;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_11_line_5 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4146 & _GEN_3981) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_11_line_5 <= _GEN_2946;
        end else begin
          cache_11_line_5 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_11_line_5 <= _GEN_2251;
      end
    end else begin
      cache_11_line_5 <= _GEN_2251;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_11_line_6 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4146 & _GEN_3983) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_11_line_6 <= _GEN_2946;
        end else begin
          cache_11_line_6 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_11_line_6 <= _GEN_2315;
      end
    end else begin
      cache_11_line_6 <= _GEN_2315;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_11_line_7 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4146 & _GEN_3985) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_11_line_7 <= _GEN_2946;
        end else begin
          cache_11_line_7 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_11_line_7 <= _GEN_2379;
      end
    end else begin
      cache_11_line_7 <= _GEN_2379;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_12_validBit <= 1'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      cache_12_validBit <= _GEN_1164;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_12_tag <= 5'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      if (6'hc == cacheLine) begin // @[Cache.scala 50:26]
        cache_12_tag <= tag; // @[Cache.scala 50:26]
      end
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_12_line_0 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4162 & _GEN_3987) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_12_line_0 <= _GEN_2946;
        end else begin
          cache_12_line_0 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_12_line_0 <= _GEN_1932;
      end
    end else begin
      cache_12_line_0 <= _GEN_1932;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_12_line_1 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4162 & _GEN_3973) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_12_line_1 <= _GEN_2946;
        end else begin
          cache_12_line_1 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_12_line_1 <= _GEN_1996;
      end
    end else begin
      cache_12_line_1 <= _GEN_1996;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_12_line_2 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4162 & _GEN_3975) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_12_line_2 <= _GEN_2946;
        end else begin
          cache_12_line_2 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_12_line_2 <= _GEN_2060;
      end
    end else begin
      cache_12_line_2 <= _GEN_2060;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_12_line_3 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4162 & _GEN_3977) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_12_line_3 <= _GEN_2946;
        end else begin
          cache_12_line_3 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_12_line_3 <= _GEN_2124;
      end
    end else begin
      cache_12_line_3 <= _GEN_2124;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_12_line_4 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4162 & _GEN_3979) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_12_line_4 <= _GEN_2946;
        end else begin
          cache_12_line_4 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_12_line_4 <= _GEN_2188;
      end
    end else begin
      cache_12_line_4 <= _GEN_2188;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_12_line_5 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4162 & _GEN_3981) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_12_line_5 <= _GEN_2946;
        end else begin
          cache_12_line_5 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_12_line_5 <= _GEN_2252;
      end
    end else begin
      cache_12_line_5 <= _GEN_2252;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_12_line_6 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4162 & _GEN_3983) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_12_line_6 <= _GEN_2946;
        end else begin
          cache_12_line_6 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_12_line_6 <= _GEN_2316;
      end
    end else begin
      cache_12_line_6 <= _GEN_2316;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_12_line_7 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4162 & _GEN_3985) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_12_line_7 <= _GEN_2946;
        end else begin
          cache_12_line_7 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_12_line_7 <= _GEN_2380;
      end
    end else begin
      cache_12_line_7 <= _GEN_2380;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_13_validBit <= 1'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      cache_13_validBit <= _GEN_1165;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_13_tag <= 5'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      if (6'hd == cacheLine) begin // @[Cache.scala 50:26]
        cache_13_tag <= tag; // @[Cache.scala 50:26]
      end
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_13_line_0 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4178 & _GEN_3987) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_13_line_0 <= _GEN_2946;
        end else begin
          cache_13_line_0 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_13_line_0 <= _GEN_1933;
      end
    end else begin
      cache_13_line_0 <= _GEN_1933;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_13_line_1 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4178 & _GEN_3973) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_13_line_1 <= _GEN_2946;
        end else begin
          cache_13_line_1 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_13_line_1 <= _GEN_1997;
      end
    end else begin
      cache_13_line_1 <= _GEN_1997;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_13_line_2 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4178 & _GEN_3975) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_13_line_2 <= _GEN_2946;
        end else begin
          cache_13_line_2 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_13_line_2 <= _GEN_2061;
      end
    end else begin
      cache_13_line_2 <= _GEN_2061;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_13_line_3 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4178 & _GEN_3977) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_13_line_3 <= _GEN_2946;
        end else begin
          cache_13_line_3 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_13_line_3 <= _GEN_2125;
      end
    end else begin
      cache_13_line_3 <= _GEN_2125;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_13_line_4 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4178 & _GEN_3979) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_13_line_4 <= _GEN_2946;
        end else begin
          cache_13_line_4 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_13_line_4 <= _GEN_2189;
      end
    end else begin
      cache_13_line_4 <= _GEN_2189;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_13_line_5 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4178 & _GEN_3981) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_13_line_5 <= _GEN_2946;
        end else begin
          cache_13_line_5 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_13_line_5 <= _GEN_2253;
      end
    end else begin
      cache_13_line_5 <= _GEN_2253;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_13_line_6 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4178 & _GEN_3983) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_13_line_6 <= _GEN_2946;
        end else begin
          cache_13_line_6 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_13_line_6 <= _GEN_2317;
      end
    end else begin
      cache_13_line_6 <= _GEN_2317;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_13_line_7 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4178 & _GEN_3985) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_13_line_7 <= _GEN_2946;
        end else begin
          cache_13_line_7 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_13_line_7 <= _GEN_2381;
      end
    end else begin
      cache_13_line_7 <= _GEN_2381;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_14_validBit <= 1'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      cache_14_validBit <= _GEN_1166;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_14_tag <= 5'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      if (6'he == cacheLine) begin // @[Cache.scala 50:26]
        cache_14_tag <= tag; // @[Cache.scala 50:26]
      end
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_14_line_0 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4194 & _GEN_3987) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_14_line_0 <= _GEN_2946;
        end else begin
          cache_14_line_0 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_14_line_0 <= _GEN_1934;
      end
    end else begin
      cache_14_line_0 <= _GEN_1934;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_14_line_1 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4194 & _GEN_3973) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_14_line_1 <= _GEN_2946;
        end else begin
          cache_14_line_1 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_14_line_1 <= _GEN_1998;
      end
    end else begin
      cache_14_line_1 <= _GEN_1998;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_14_line_2 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4194 & _GEN_3975) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_14_line_2 <= _GEN_2946;
        end else begin
          cache_14_line_2 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_14_line_2 <= _GEN_2062;
      end
    end else begin
      cache_14_line_2 <= _GEN_2062;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_14_line_3 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4194 & _GEN_3977) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_14_line_3 <= _GEN_2946;
        end else begin
          cache_14_line_3 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_14_line_3 <= _GEN_2126;
      end
    end else begin
      cache_14_line_3 <= _GEN_2126;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_14_line_4 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4194 & _GEN_3979) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_14_line_4 <= _GEN_2946;
        end else begin
          cache_14_line_4 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_14_line_4 <= _GEN_2190;
      end
    end else begin
      cache_14_line_4 <= _GEN_2190;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_14_line_5 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4194 & _GEN_3981) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_14_line_5 <= _GEN_2946;
        end else begin
          cache_14_line_5 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_14_line_5 <= _GEN_2254;
      end
    end else begin
      cache_14_line_5 <= _GEN_2254;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_14_line_6 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4194 & _GEN_3983) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_14_line_6 <= _GEN_2946;
        end else begin
          cache_14_line_6 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_14_line_6 <= _GEN_2318;
      end
    end else begin
      cache_14_line_6 <= _GEN_2318;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_14_line_7 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4194 & _GEN_3985) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_14_line_7 <= _GEN_2946;
        end else begin
          cache_14_line_7 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_14_line_7 <= _GEN_2382;
      end
    end else begin
      cache_14_line_7 <= _GEN_2382;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_15_validBit <= 1'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      cache_15_validBit <= _GEN_1167;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_15_tag <= 5'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      if (6'hf == cacheLine) begin // @[Cache.scala 50:26]
        cache_15_tag <= tag; // @[Cache.scala 50:26]
      end
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_15_line_0 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4210 & _GEN_3987) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_15_line_0 <= _GEN_2946;
        end else begin
          cache_15_line_0 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_15_line_0 <= _GEN_1935;
      end
    end else begin
      cache_15_line_0 <= _GEN_1935;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_15_line_1 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4210 & _GEN_3973) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_15_line_1 <= _GEN_2946;
        end else begin
          cache_15_line_1 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_15_line_1 <= _GEN_1999;
      end
    end else begin
      cache_15_line_1 <= _GEN_1999;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_15_line_2 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4210 & _GEN_3975) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_15_line_2 <= _GEN_2946;
        end else begin
          cache_15_line_2 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_15_line_2 <= _GEN_2063;
      end
    end else begin
      cache_15_line_2 <= _GEN_2063;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_15_line_3 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4210 & _GEN_3977) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_15_line_3 <= _GEN_2946;
        end else begin
          cache_15_line_3 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_15_line_3 <= _GEN_2127;
      end
    end else begin
      cache_15_line_3 <= _GEN_2127;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_15_line_4 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4210 & _GEN_3979) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_15_line_4 <= _GEN_2946;
        end else begin
          cache_15_line_4 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_15_line_4 <= _GEN_2191;
      end
    end else begin
      cache_15_line_4 <= _GEN_2191;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_15_line_5 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4210 & _GEN_3981) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_15_line_5 <= _GEN_2946;
        end else begin
          cache_15_line_5 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_15_line_5 <= _GEN_2255;
      end
    end else begin
      cache_15_line_5 <= _GEN_2255;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_15_line_6 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4210 & _GEN_3983) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_15_line_6 <= _GEN_2946;
        end else begin
          cache_15_line_6 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_15_line_6 <= _GEN_2319;
      end
    end else begin
      cache_15_line_6 <= _GEN_2319;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_15_line_7 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4210 & _GEN_3985) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_15_line_7 <= _GEN_2946;
        end else begin
          cache_15_line_7 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_15_line_7 <= _GEN_2383;
      end
    end else begin
      cache_15_line_7 <= _GEN_2383;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_16_validBit <= 1'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      cache_16_validBit <= _GEN_1168;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_16_tag <= 5'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      if (6'h10 == cacheLine) begin // @[Cache.scala 50:26]
        cache_16_tag <= tag; // @[Cache.scala 50:26]
      end
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_16_line_0 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4226 & _GEN_3987) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_16_line_0 <= _GEN_2946;
        end else begin
          cache_16_line_0 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_16_line_0 <= _GEN_1936;
      end
    end else begin
      cache_16_line_0 <= _GEN_1936;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_16_line_1 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4226 & _GEN_3973) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_16_line_1 <= _GEN_2946;
        end else begin
          cache_16_line_1 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_16_line_1 <= _GEN_2000;
      end
    end else begin
      cache_16_line_1 <= _GEN_2000;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_16_line_2 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4226 & _GEN_3975) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_16_line_2 <= _GEN_2946;
        end else begin
          cache_16_line_2 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_16_line_2 <= _GEN_2064;
      end
    end else begin
      cache_16_line_2 <= _GEN_2064;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_16_line_3 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4226 & _GEN_3977) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_16_line_3 <= _GEN_2946;
        end else begin
          cache_16_line_3 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_16_line_3 <= _GEN_2128;
      end
    end else begin
      cache_16_line_3 <= _GEN_2128;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_16_line_4 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4226 & _GEN_3979) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_16_line_4 <= _GEN_2946;
        end else begin
          cache_16_line_4 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_16_line_4 <= _GEN_2192;
      end
    end else begin
      cache_16_line_4 <= _GEN_2192;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_16_line_5 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4226 & _GEN_3981) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_16_line_5 <= _GEN_2946;
        end else begin
          cache_16_line_5 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_16_line_5 <= _GEN_2256;
      end
    end else begin
      cache_16_line_5 <= _GEN_2256;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_16_line_6 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4226 & _GEN_3983) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_16_line_6 <= _GEN_2946;
        end else begin
          cache_16_line_6 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_16_line_6 <= _GEN_2320;
      end
    end else begin
      cache_16_line_6 <= _GEN_2320;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_16_line_7 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4226 & _GEN_3985) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_16_line_7 <= _GEN_2946;
        end else begin
          cache_16_line_7 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_16_line_7 <= _GEN_2384;
      end
    end else begin
      cache_16_line_7 <= _GEN_2384;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_17_validBit <= 1'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      cache_17_validBit <= _GEN_1169;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_17_tag <= 5'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      if (6'h11 == cacheLine) begin // @[Cache.scala 50:26]
        cache_17_tag <= tag; // @[Cache.scala 50:26]
      end
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_17_line_0 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4242 & _GEN_3987) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_17_line_0 <= _GEN_2946;
        end else begin
          cache_17_line_0 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_17_line_0 <= _GEN_1937;
      end
    end else begin
      cache_17_line_0 <= _GEN_1937;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_17_line_1 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4242 & _GEN_3973) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_17_line_1 <= _GEN_2946;
        end else begin
          cache_17_line_1 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_17_line_1 <= _GEN_2001;
      end
    end else begin
      cache_17_line_1 <= _GEN_2001;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_17_line_2 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4242 & _GEN_3975) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_17_line_2 <= _GEN_2946;
        end else begin
          cache_17_line_2 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_17_line_2 <= _GEN_2065;
      end
    end else begin
      cache_17_line_2 <= _GEN_2065;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_17_line_3 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4242 & _GEN_3977) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_17_line_3 <= _GEN_2946;
        end else begin
          cache_17_line_3 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_17_line_3 <= _GEN_2129;
      end
    end else begin
      cache_17_line_3 <= _GEN_2129;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_17_line_4 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4242 & _GEN_3979) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_17_line_4 <= _GEN_2946;
        end else begin
          cache_17_line_4 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_17_line_4 <= _GEN_2193;
      end
    end else begin
      cache_17_line_4 <= _GEN_2193;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_17_line_5 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4242 & _GEN_3981) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_17_line_5 <= _GEN_2946;
        end else begin
          cache_17_line_5 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_17_line_5 <= _GEN_2257;
      end
    end else begin
      cache_17_line_5 <= _GEN_2257;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_17_line_6 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4242 & _GEN_3983) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_17_line_6 <= _GEN_2946;
        end else begin
          cache_17_line_6 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_17_line_6 <= _GEN_2321;
      end
    end else begin
      cache_17_line_6 <= _GEN_2321;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_17_line_7 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4242 & _GEN_3985) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_17_line_7 <= _GEN_2946;
        end else begin
          cache_17_line_7 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_17_line_7 <= _GEN_2385;
      end
    end else begin
      cache_17_line_7 <= _GEN_2385;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_18_validBit <= 1'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      cache_18_validBit <= _GEN_1170;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_18_tag <= 5'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      if (6'h12 == cacheLine) begin // @[Cache.scala 50:26]
        cache_18_tag <= tag; // @[Cache.scala 50:26]
      end
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_18_line_0 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4258 & _GEN_3987) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_18_line_0 <= _GEN_2946;
        end else begin
          cache_18_line_0 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_18_line_0 <= _GEN_1938;
      end
    end else begin
      cache_18_line_0 <= _GEN_1938;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_18_line_1 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4258 & _GEN_3973) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_18_line_1 <= _GEN_2946;
        end else begin
          cache_18_line_1 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_18_line_1 <= _GEN_2002;
      end
    end else begin
      cache_18_line_1 <= _GEN_2002;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_18_line_2 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4258 & _GEN_3975) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_18_line_2 <= _GEN_2946;
        end else begin
          cache_18_line_2 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_18_line_2 <= _GEN_2066;
      end
    end else begin
      cache_18_line_2 <= _GEN_2066;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_18_line_3 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4258 & _GEN_3977) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_18_line_3 <= _GEN_2946;
        end else begin
          cache_18_line_3 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_18_line_3 <= _GEN_2130;
      end
    end else begin
      cache_18_line_3 <= _GEN_2130;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_18_line_4 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4258 & _GEN_3979) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_18_line_4 <= _GEN_2946;
        end else begin
          cache_18_line_4 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_18_line_4 <= _GEN_2194;
      end
    end else begin
      cache_18_line_4 <= _GEN_2194;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_18_line_5 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4258 & _GEN_3981) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_18_line_5 <= _GEN_2946;
        end else begin
          cache_18_line_5 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_18_line_5 <= _GEN_2258;
      end
    end else begin
      cache_18_line_5 <= _GEN_2258;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_18_line_6 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4258 & _GEN_3983) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_18_line_6 <= _GEN_2946;
        end else begin
          cache_18_line_6 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_18_line_6 <= _GEN_2322;
      end
    end else begin
      cache_18_line_6 <= _GEN_2322;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_18_line_7 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4258 & _GEN_3985) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_18_line_7 <= _GEN_2946;
        end else begin
          cache_18_line_7 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_18_line_7 <= _GEN_2386;
      end
    end else begin
      cache_18_line_7 <= _GEN_2386;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_19_validBit <= 1'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      cache_19_validBit <= _GEN_1171;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_19_tag <= 5'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      if (6'h13 == cacheLine) begin // @[Cache.scala 50:26]
        cache_19_tag <= tag; // @[Cache.scala 50:26]
      end
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_19_line_0 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4274 & _GEN_3987) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_19_line_0 <= _GEN_2946;
        end else begin
          cache_19_line_0 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_19_line_0 <= _GEN_1939;
      end
    end else begin
      cache_19_line_0 <= _GEN_1939;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_19_line_1 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4274 & _GEN_3973) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_19_line_1 <= _GEN_2946;
        end else begin
          cache_19_line_1 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_19_line_1 <= _GEN_2003;
      end
    end else begin
      cache_19_line_1 <= _GEN_2003;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_19_line_2 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4274 & _GEN_3975) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_19_line_2 <= _GEN_2946;
        end else begin
          cache_19_line_2 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_19_line_2 <= _GEN_2067;
      end
    end else begin
      cache_19_line_2 <= _GEN_2067;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_19_line_3 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4274 & _GEN_3977) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_19_line_3 <= _GEN_2946;
        end else begin
          cache_19_line_3 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_19_line_3 <= _GEN_2131;
      end
    end else begin
      cache_19_line_3 <= _GEN_2131;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_19_line_4 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4274 & _GEN_3979) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_19_line_4 <= _GEN_2946;
        end else begin
          cache_19_line_4 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_19_line_4 <= _GEN_2195;
      end
    end else begin
      cache_19_line_4 <= _GEN_2195;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_19_line_5 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4274 & _GEN_3981) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_19_line_5 <= _GEN_2946;
        end else begin
          cache_19_line_5 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_19_line_5 <= _GEN_2259;
      end
    end else begin
      cache_19_line_5 <= _GEN_2259;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_19_line_6 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4274 & _GEN_3983) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_19_line_6 <= _GEN_2946;
        end else begin
          cache_19_line_6 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_19_line_6 <= _GEN_2323;
      end
    end else begin
      cache_19_line_6 <= _GEN_2323;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_19_line_7 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4274 & _GEN_3985) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_19_line_7 <= _GEN_2946;
        end else begin
          cache_19_line_7 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_19_line_7 <= _GEN_2387;
      end
    end else begin
      cache_19_line_7 <= _GEN_2387;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_20_validBit <= 1'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      cache_20_validBit <= _GEN_1172;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_20_tag <= 5'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      if (6'h14 == cacheLine) begin // @[Cache.scala 50:26]
        cache_20_tag <= tag; // @[Cache.scala 50:26]
      end
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_20_line_0 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4290 & _GEN_3987) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_20_line_0 <= _GEN_2946;
        end else begin
          cache_20_line_0 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_20_line_0 <= _GEN_1940;
      end
    end else begin
      cache_20_line_0 <= _GEN_1940;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_20_line_1 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4290 & _GEN_3973) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_20_line_1 <= _GEN_2946;
        end else begin
          cache_20_line_1 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_20_line_1 <= _GEN_2004;
      end
    end else begin
      cache_20_line_1 <= _GEN_2004;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_20_line_2 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4290 & _GEN_3975) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_20_line_2 <= _GEN_2946;
        end else begin
          cache_20_line_2 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_20_line_2 <= _GEN_2068;
      end
    end else begin
      cache_20_line_2 <= _GEN_2068;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_20_line_3 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4290 & _GEN_3977) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_20_line_3 <= _GEN_2946;
        end else begin
          cache_20_line_3 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_20_line_3 <= _GEN_2132;
      end
    end else begin
      cache_20_line_3 <= _GEN_2132;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_20_line_4 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4290 & _GEN_3979) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_20_line_4 <= _GEN_2946;
        end else begin
          cache_20_line_4 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_20_line_4 <= _GEN_2196;
      end
    end else begin
      cache_20_line_4 <= _GEN_2196;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_20_line_5 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4290 & _GEN_3981) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_20_line_5 <= _GEN_2946;
        end else begin
          cache_20_line_5 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_20_line_5 <= _GEN_2260;
      end
    end else begin
      cache_20_line_5 <= _GEN_2260;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_20_line_6 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4290 & _GEN_3983) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_20_line_6 <= _GEN_2946;
        end else begin
          cache_20_line_6 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_20_line_6 <= _GEN_2324;
      end
    end else begin
      cache_20_line_6 <= _GEN_2324;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_20_line_7 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4290 & _GEN_3985) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_20_line_7 <= _GEN_2946;
        end else begin
          cache_20_line_7 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_20_line_7 <= _GEN_2388;
      end
    end else begin
      cache_20_line_7 <= _GEN_2388;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_21_validBit <= 1'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      cache_21_validBit <= _GEN_1173;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_21_tag <= 5'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      if (6'h15 == cacheLine) begin // @[Cache.scala 50:26]
        cache_21_tag <= tag; // @[Cache.scala 50:26]
      end
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_21_line_0 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4306 & _GEN_3987) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_21_line_0 <= _GEN_2946;
        end else begin
          cache_21_line_0 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_21_line_0 <= _GEN_1941;
      end
    end else begin
      cache_21_line_0 <= _GEN_1941;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_21_line_1 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4306 & _GEN_3973) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_21_line_1 <= _GEN_2946;
        end else begin
          cache_21_line_1 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_21_line_1 <= _GEN_2005;
      end
    end else begin
      cache_21_line_1 <= _GEN_2005;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_21_line_2 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4306 & _GEN_3975) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_21_line_2 <= _GEN_2946;
        end else begin
          cache_21_line_2 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_21_line_2 <= _GEN_2069;
      end
    end else begin
      cache_21_line_2 <= _GEN_2069;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_21_line_3 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4306 & _GEN_3977) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_21_line_3 <= _GEN_2946;
        end else begin
          cache_21_line_3 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_21_line_3 <= _GEN_2133;
      end
    end else begin
      cache_21_line_3 <= _GEN_2133;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_21_line_4 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4306 & _GEN_3979) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_21_line_4 <= _GEN_2946;
        end else begin
          cache_21_line_4 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_21_line_4 <= _GEN_2197;
      end
    end else begin
      cache_21_line_4 <= _GEN_2197;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_21_line_5 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4306 & _GEN_3981) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_21_line_5 <= _GEN_2946;
        end else begin
          cache_21_line_5 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_21_line_5 <= _GEN_2261;
      end
    end else begin
      cache_21_line_5 <= _GEN_2261;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_21_line_6 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4306 & _GEN_3983) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_21_line_6 <= _GEN_2946;
        end else begin
          cache_21_line_6 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_21_line_6 <= _GEN_2325;
      end
    end else begin
      cache_21_line_6 <= _GEN_2325;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_21_line_7 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4306 & _GEN_3985) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_21_line_7 <= _GEN_2946;
        end else begin
          cache_21_line_7 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_21_line_7 <= _GEN_2389;
      end
    end else begin
      cache_21_line_7 <= _GEN_2389;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_22_validBit <= 1'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      cache_22_validBit <= _GEN_1174;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_22_tag <= 5'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      if (6'h16 == cacheLine) begin // @[Cache.scala 50:26]
        cache_22_tag <= tag; // @[Cache.scala 50:26]
      end
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_22_line_0 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4322 & _GEN_3987) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_22_line_0 <= _GEN_2946;
        end else begin
          cache_22_line_0 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_22_line_0 <= _GEN_1942;
      end
    end else begin
      cache_22_line_0 <= _GEN_1942;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_22_line_1 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4322 & _GEN_3973) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_22_line_1 <= _GEN_2946;
        end else begin
          cache_22_line_1 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_22_line_1 <= _GEN_2006;
      end
    end else begin
      cache_22_line_1 <= _GEN_2006;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_22_line_2 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4322 & _GEN_3975) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_22_line_2 <= _GEN_2946;
        end else begin
          cache_22_line_2 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_22_line_2 <= _GEN_2070;
      end
    end else begin
      cache_22_line_2 <= _GEN_2070;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_22_line_3 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4322 & _GEN_3977) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_22_line_3 <= _GEN_2946;
        end else begin
          cache_22_line_3 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_22_line_3 <= _GEN_2134;
      end
    end else begin
      cache_22_line_3 <= _GEN_2134;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_22_line_4 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4322 & _GEN_3979) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_22_line_4 <= _GEN_2946;
        end else begin
          cache_22_line_4 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_22_line_4 <= _GEN_2198;
      end
    end else begin
      cache_22_line_4 <= _GEN_2198;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_22_line_5 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4322 & _GEN_3981) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_22_line_5 <= _GEN_2946;
        end else begin
          cache_22_line_5 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_22_line_5 <= _GEN_2262;
      end
    end else begin
      cache_22_line_5 <= _GEN_2262;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_22_line_6 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4322 & _GEN_3983) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_22_line_6 <= _GEN_2946;
        end else begin
          cache_22_line_6 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_22_line_6 <= _GEN_2326;
      end
    end else begin
      cache_22_line_6 <= _GEN_2326;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_22_line_7 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4322 & _GEN_3985) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_22_line_7 <= _GEN_2946;
        end else begin
          cache_22_line_7 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_22_line_7 <= _GEN_2390;
      end
    end else begin
      cache_22_line_7 <= _GEN_2390;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_23_validBit <= 1'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      cache_23_validBit <= _GEN_1175;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_23_tag <= 5'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      if (6'h17 == cacheLine) begin // @[Cache.scala 50:26]
        cache_23_tag <= tag; // @[Cache.scala 50:26]
      end
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_23_line_0 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4338 & _GEN_3987) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_23_line_0 <= _GEN_2946;
        end else begin
          cache_23_line_0 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_23_line_0 <= _GEN_1943;
      end
    end else begin
      cache_23_line_0 <= _GEN_1943;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_23_line_1 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4338 & _GEN_3973) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_23_line_1 <= _GEN_2946;
        end else begin
          cache_23_line_1 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_23_line_1 <= _GEN_2007;
      end
    end else begin
      cache_23_line_1 <= _GEN_2007;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_23_line_2 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4338 & _GEN_3975) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_23_line_2 <= _GEN_2946;
        end else begin
          cache_23_line_2 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_23_line_2 <= _GEN_2071;
      end
    end else begin
      cache_23_line_2 <= _GEN_2071;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_23_line_3 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4338 & _GEN_3977) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_23_line_3 <= _GEN_2946;
        end else begin
          cache_23_line_3 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_23_line_3 <= _GEN_2135;
      end
    end else begin
      cache_23_line_3 <= _GEN_2135;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_23_line_4 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4338 & _GEN_3979) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_23_line_4 <= _GEN_2946;
        end else begin
          cache_23_line_4 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_23_line_4 <= _GEN_2199;
      end
    end else begin
      cache_23_line_4 <= _GEN_2199;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_23_line_5 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4338 & _GEN_3981) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_23_line_5 <= _GEN_2946;
        end else begin
          cache_23_line_5 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_23_line_5 <= _GEN_2263;
      end
    end else begin
      cache_23_line_5 <= _GEN_2263;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_23_line_6 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4338 & _GEN_3983) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_23_line_6 <= _GEN_2946;
        end else begin
          cache_23_line_6 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_23_line_6 <= _GEN_2327;
      end
    end else begin
      cache_23_line_6 <= _GEN_2327;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_23_line_7 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4338 & _GEN_3985) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_23_line_7 <= _GEN_2946;
        end else begin
          cache_23_line_7 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_23_line_7 <= _GEN_2391;
      end
    end else begin
      cache_23_line_7 <= _GEN_2391;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_24_validBit <= 1'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      cache_24_validBit <= _GEN_1176;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_24_tag <= 5'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      if (6'h18 == cacheLine) begin // @[Cache.scala 50:26]
        cache_24_tag <= tag; // @[Cache.scala 50:26]
      end
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_24_line_0 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4354 & _GEN_3987) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_24_line_0 <= _GEN_2946;
        end else begin
          cache_24_line_0 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_24_line_0 <= _GEN_1944;
      end
    end else begin
      cache_24_line_0 <= _GEN_1944;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_24_line_1 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4354 & _GEN_3973) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_24_line_1 <= _GEN_2946;
        end else begin
          cache_24_line_1 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_24_line_1 <= _GEN_2008;
      end
    end else begin
      cache_24_line_1 <= _GEN_2008;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_24_line_2 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4354 & _GEN_3975) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_24_line_2 <= _GEN_2946;
        end else begin
          cache_24_line_2 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_24_line_2 <= _GEN_2072;
      end
    end else begin
      cache_24_line_2 <= _GEN_2072;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_24_line_3 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4354 & _GEN_3977) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_24_line_3 <= _GEN_2946;
        end else begin
          cache_24_line_3 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_24_line_3 <= _GEN_2136;
      end
    end else begin
      cache_24_line_3 <= _GEN_2136;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_24_line_4 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4354 & _GEN_3979) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_24_line_4 <= _GEN_2946;
        end else begin
          cache_24_line_4 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_24_line_4 <= _GEN_2200;
      end
    end else begin
      cache_24_line_4 <= _GEN_2200;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_24_line_5 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4354 & _GEN_3981) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_24_line_5 <= _GEN_2946;
        end else begin
          cache_24_line_5 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_24_line_5 <= _GEN_2264;
      end
    end else begin
      cache_24_line_5 <= _GEN_2264;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_24_line_6 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4354 & _GEN_3983) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_24_line_6 <= _GEN_2946;
        end else begin
          cache_24_line_6 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_24_line_6 <= _GEN_2328;
      end
    end else begin
      cache_24_line_6 <= _GEN_2328;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_24_line_7 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4354 & _GEN_3985) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_24_line_7 <= _GEN_2946;
        end else begin
          cache_24_line_7 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_24_line_7 <= _GEN_2392;
      end
    end else begin
      cache_24_line_7 <= _GEN_2392;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_25_validBit <= 1'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      cache_25_validBit <= _GEN_1177;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_25_tag <= 5'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      if (6'h19 == cacheLine) begin // @[Cache.scala 50:26]
        cache_25_tag <= tag; // @[Cache.scala 50:26]
      end
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_25_line_0 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4370 & _GEN_3987) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_25_line_0 <= _GEN_2946;
        end else begin
          cache_25_line_0 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_25_line_0 <= _GEN_1945;
      end
    end else begin
      cache_25_line_0 <= _GEN_1945;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_25_line_1 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4370 & _GEN_3973) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_25_line_1 <= _GEN_2946;
        end else begin
          cache_25_line_1 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_25_line_1 <= _GEN_2009;
      end
    end else begin
      cache_25_line_1 <= _GEN_2009;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_25_line_2 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4370 & _GEN_3975) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_25_line_2 <= _GEN_2946;
        end else begin
          cache_25_line_2 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_25_line_2 <= _GEN_2073;
      end
    end else begin
      cache_25_line_2 <= _GEN_2073;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_25_line_3 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4370 & _GEN_3977) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_25_line_3 <= _GEN_2946;
        end else begin
          cache_25_line_3 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_25_line_3 <= _GEN_2137;
      end
    end else begin
      cache_25_line_3 <= _GEN_2137;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_25_line_4 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4370 & _GEN_3979) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_25_line_4 <= _GEN_2946;
        end else begin
          cache_25_line_4 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_25_line_4 <= _GEN_2201;
      end
    end else begin
      cache_25_line_4 <= _GEN_2201;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_25_line_5 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4370 & _GEN_3981) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_25_line_5 <= _GEN_2946;
        end else begin
          cache_25_line_5 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_25_line_5 <= _GEN_2265;
      end
    end else begin
      cache_25_line_5 <= _GEN_2265;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_25_line_6 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4370 & _GEN_3983) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_25_line_6 <= _GEN_2946;
        end else begin
          cache_25_line_6 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_25_line_6 <= _GEN_2329;
      end
    end else begin
      cache_25_line_6 <= _GEN_2329;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_25_line_7 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4370 & _GEN_3985) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_25_line_7 <= _GEN_2946;
        end else begin
          cache_25_line_7 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_25_line_7 <= _GEN_2393;
      end
    end else begin
      cache_25_line_7 <= _GEN_2393;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_26_validBit <= 1'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      cache_26_validBit <= _GEN_1178;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_26_tag <= 5'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      if (6'h1a == cacheLine) begin // @[Cache.scala 50:26]
        cache_26_tag <= tag; // @[Cache.scala 50:26]
      end
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_26_line_0 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4386 & _GEN_3987) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_26_line_0 <= _GEN_2946;
        end else begin
          cache_26_line_0 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_26_line_0 <= _GEN_1946;
      end
    end else begin
      cache_26_line_0 <= _GEN_1946;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_26_line_1 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4386 & _GEN_3973) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_26_line_1 <= _GEN_2946;
        end else begin
          cache_26_line_1 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_26_line_1 <= _GEN_2010;
      end
    end else begin
      cache_26_line_1 <= _GEN_2010;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_26_line_2 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4386 & _GEN_3975) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_26_line_2 <= _GEN_2946;
        end else begin
          cache_26_line_2 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_26_line_2 <= _GEN_2074;
      end
    end else begin
      cache_26_line_2 <= _GEN_2074;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_26_line_3 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4386 & _GEN_3977) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_26_line_3 <= _GEN_2946;
        end else begin
          cache_26_line_3 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_26_line_3 <= _GEN_2138;
      end
    end else begin
      cache_26_line_3 <= _GEN_2138;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_26_line_4 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4386 & _GEN_3979) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_26_line_4 <= _GEN_2946;
        end else begin
          cache_26_line_4 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_26_line_4 <= _GEN_2202;
      end
    end else begin
      cache_26_line_4 <= _GEN_2202;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_26_line_5 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4386 & _GEN_3981) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_26_line_5 <= _GEN_2946;
        end else begin
          cache_26_line_5 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_26_line_5 <= _GEN_2266;
      end
    end else begin
      cache_26_line_5 <= _GEN_2266;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_26_line_6 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4386 & _GEN_3983) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_26_line_6 <= _GEN_2946;
        end else begin
          cache_26_line_6 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_26_line_6 <= _GEN_2330;
      end
    end else begin
      cache_26_line_6 <= _GEN_2330;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_26_line_7 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4386 & _GEN_3985) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_26_line_7 <= _GEN_2946;
        end else begin
          cache_26_line_7 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_26_line_7 <= _GEN_2394;
      end
    end else begin
      cache_26_line_7 <= _GEN_2394;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_27_validBit <= 1'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      cache_27_validBit <= _GEN_1179;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_27_tag <= 5'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      if (6'h1b == cacheLine) begin // @[Cache.scala 50:26]
        cache_27_tag <= tag; // @[Cache.scala 50:26]
      end
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_27_line_0 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4402 & _GEN_3987) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_27_line_0 <= _GEN_2946;
        end else begin
          cache_27_line_0 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_27_line_0 <= _GEN_1947;
      end
    end else begin
      cache_27_line_0 <= _GEN_1947;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_27_line_1 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4402 & _GEN_3973) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_27_line_1 <= _GEN_2946;
        end else begin
          cache_27_line_1 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_27_line_1 <= _GEN_2011;
      end
    end else begin
      cache_27_line_1 <= _GEN_2011;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_27_line_2 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4402 & _GEN_3975) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_27_line_2 <= _GEN_2946;
        end else begin
          cache_27_line_2 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_27_line_2 <= _GEN_2075;
      end
    end else begin
      cache_27_line_2 <= _GEN_2075;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_27_line_3 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4402 & _GEN_3977) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_27_line_3 <= _GEN_2946;
        end else begin
          cache_27_line_3 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_27_line_3 <= _GEN_2139;
      end
    end else begin
      cache_27_line_3 <= _GEN_2139;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_27_line_4 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4402 & _GEN_3979) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_27_line_4 <= _GEN_2946;
        end else begin
          cache_27_line_4 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_27_line_4 <= _GEN_2203;
      end
    end else begin
      cache_27_line_4 <= _GEN_2203;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_27_line_5 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4402 & _GEN_3981) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_27_line_5 <= _GEN_2946;
        end else begin
          cache_27_line_5 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_27_line_5 <= _GEN_2267;
      end
    end else begin
      cache_27_line_5 <= _GEN_2267;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_27_line_6 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4402 & _GEN_3983) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_27_line_6 <= _GEN_2946;
        end else begin
          cache_27_line_6 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_27_line_6 <= _GEN_2331;
      end
    end else begin
      cache_27_line_6 <= _GEN_2331;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_27_line_7 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4402 & _GEN_3985) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_27_line_7 <= _GEN_2946;
        end else begin
          cache_27_line_7 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_27_line_7 <= _GEN_2395;
      end
    end else begin
      cache_27_line_7 <= _GEN_2395;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_28_validBit <= 1'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      cache_28_validBit <= _GEN_1180;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_28_tag <= 5'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      if (6'h1c == cacheLine) begin // @[Cache.scala 50:26]
        cache_28_tag <= tag; // @[Cache.scala 50:26]
      end
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_28_line_0 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4418 & _GEN_3987) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_28_line_0 <= _GEN_2946;
        end else begin
          cache_28_line_0 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_28_line_0 <= _GEN_1948;
      end
    end else begin
      cache_28_line_0 <= _GEN_1948;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_28_line_1 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4418 & _GEN_3973) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_28_line_1 <= _GEN_2946;
        end else begin
          cache_28_line_1 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_28_line_1 <= _GEN_2012;
      end
    end else begin
      cache_28_line_1 <= _GEN_2012;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_28_line_2 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4418 & _GEN_3975) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_28_line_2 <= _GEN_2946;
        end else begin
          cache_28_line_2 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_28_line_2 <= _GEN_2076;
      end
    end else begin
      cache_28_line_2 <= _GEN_2076;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_28_line_3 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4418 & _GEN_3977) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_28_line_3 <= _GEN_2946;
        end else begin
          cache_28_line_3 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_28_line_3 <= _GEN_2140;
      end
    end else begin
      cache_28_line_3 <= _GEN_2140;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_28_line_4 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4418 & _GEN_3979) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_28_line_4 <= _GEN_2946;
        end else begin
          cache_28_line_4 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_28_line_4 <= _GEN_2204;
      end
    end else begin
      cache_28_line_4 <= _GEN_2204;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_28_line_5 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4418 & _GEN_3981) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_28_line_5 <= _GEN_2946;
        end else begin
          cache_28_line_5 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_28_line_5 <= _GEN_2268;
      end
    end else begin
      cache_28_line_5 <= _GEN_2268;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_28_line_6 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4418 & _GEN_3983) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_28_line_6 <= _GEN_2946;
        end else begin
          cache_28_line_6 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_28_line_6 <= _GEN_2332;
      end
    end else begin
      cache_28_line_6 <= _GEN_2332;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_28_line_7 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4418 & _GEN_3985) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_28_line_7 <= _GEN_2946;
        end else begin
          cache_28_line_7 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_28_line_7 <= _GEN_2396;
      end
    end else begin
      cache_28_line_7 <= _GEN_2396;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_29_validBit <= 1'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      cache_29_validBit <= _GEN_1181;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_29_tag <= 5'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      if (6'h1d == cacheLine) begin // @[Cache.scala 50:26]
        cache_29_tag <= tag; // @[Cache.scala 50:26]
      end
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_29_line_0 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4434 & _GEN_3987) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_29_line_0 <= _GEN_2946;
        end else begin
          cache_29_line_0 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_29_line_0 <= _GEN_1949;
      end
    end else begin
      cache_29_line_0 <= _GEN_1949;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_29_line_1 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4434 & _GEN_3973) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_29_line_1 <= _GEN_2946;
        end else begin
          cache_29_line_1 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_29_line_1 <= _GEN_2013;
      end
    end else begin
      cache_29_line_1 <= _GEN_2013;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_29_line_2 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4434 & _GEN_3975) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_29_line_2 <= _GEN_2946;
        end else begin
          cache_29_line_2 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_29_line_2 <= _GEN_2077;
      end
    end else begin
      cache_29_line_2 <= _GEN_2077;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_29_line_3 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4434 & _GEN_3977) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_29_line_3 <= _GEN_2946;
        end else begin
          cache_29_line_3 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_29_line_3 <= _GEN_2141;
      end
    end else begin
      cache_29_line_3 <= _GEN_2141;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_29_line_4 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4434 & _GEN_3979) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_29_line_4 <= _GEN_2946;
        end else begin
          cache_29_line_4 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_29_line_4 <= _GEN_2205;
      end
    end else begin
      cache_29_line_4 <= _GEN_2205;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_29_line_5 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4434 & _GEN_3981) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_29_line_5 <= _GEN_2946;
        end else begin
          cache_29_line_5 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_29_line_5 <= _GEN_2269;
      end
    end else begin
      cache_29_line_5 <= _GEN_2269;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_29_line_6 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4434 & _GEN_3983) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_29_line_6 <= _GEN_2946;
        end else begin
          cache_29_line_6 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_29_line_6 <= _GEN_2333;
      end
    end else begin
      cache_29_line_6 <= _GEN_2333;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_29_line_7 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4434 & _GEN_3985) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_29_line_7 <= _GEN_2946;
        end else begin
          cache_29_line_7 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_29_line_7 <= _GEN_2397;
      end
    end else begin
      cache_29_line_7 <= _GEN_2397;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_30_validBit <= 1'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      cache_30_validBit <= _GEN_1182;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_30_tag <= 5'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      if (6'h1e == cacheLine) begin // @[Cache.scala 50:26]
        cache_30_tag <= tag; // @[Cache.scala 50:26]
      end
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_30_line_0 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4450 & _GEN_3987) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_30_line_0 <= _GEN_2946;
        end else begin
          cache_30_line_0 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_30_line_0 <= _GEN_1950;
      end
    end else begin
      cache_30_line_0 <= _GEN_1950;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_30_line_1 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4450 & _GEN_3973) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_30_line_1 <= _GEN_2946;
        end else begin
          cache_30_line_1 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_30_line_1 <= _GEN_2014;
      end
    end else begin
      cache_30_line_1 <= _GEN_2014;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_30_line_2 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4450 & _GEN_3975) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_30_line_2 <= _GEN_2946;
        end else begin
          cache_30_line_2 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_30_line_2 <= _GEN_2078;
      end
    end else begin
      cache_30_line_2 <= _GEN_2078;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_30_line_3 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4450 & _GEN_3977) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_30_line_3 <= _GEN_2946;
        end else begin
          cache_30_line_3 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_30_line_3 <= _GEN_2142;
      end
    end else begin
      cache_30_line_3 <= _GEN_2142;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_30_line_4 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4450 & _GEN_3979) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_30_line_4 <= _GEN_2946;
        end else begin
          cache_30_line_4 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_30_line_4 <= _GEN_2206;
      end
    end else begin
      cache_30_line_4 <= _GEN_2206;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_30_line_5 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4450 & _GEN_3981) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_30_line_5 <= _GEN_2946;
        end else begin
          cache_30_line_5 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_30_line_5 <= _GEN_2270;
      end
    end else begin
      cache_30_line_5 <= _GEN_2270;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_30_line_6 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4450 & _GEN_3983) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_30_line_6 <= _GEN_2946;
        end else begin
          cache_30_line_6 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_30_line_6 <= _GEN_2334;
      end
    end else begin
      cache_30_line_6 <= _GEN_2334;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_30_line_7 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4450 & _GEN_3985) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_30_line_7 <= _GEN_2946;
        end else begin
          cache_30_line_7 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_30_line_7 <= _GEN_2398;
      end
    end else begin
      cache_30_line_7 <= _GEN_2398;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_31_validBit <= 1'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      cache_31_validBit <= _GEN_1183;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_31_tag <= 5'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      if (6'h1f == cacheLine) begin // @[Cache.scala 50:26]
        cache_31_tag <= tag; // @[Cache.scala 50:26]
      end
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_31_line_0 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4466 & _GEN_3987) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_31_line_0 <= _GEN_2946;
        end else begin
          cache_31_line_0 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_31_line_0 <= _GEN_1951;
      end
    end else begin
      cache_31_line_0 <= _GEN_1951;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_31_line_1 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4466 & _GEN_3973) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_31_line_1 <= _GEN_2946;
        end else begin
          cache_31_line_1 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_31_line_1 <= _GEN_2015;
      end
    end else begin
      cache_31_line_1 <= _GEN_2015;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_31_line_2 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4466 & _GEN_3975) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_31_line_2 <= _GEN_2946;
        end else begin
          cache_31_line_2 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_31_line_2 <= _GEN_2079;
      end
    end else begin
      cache_31_line_2 <= _GEN_2079;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_31_line_3 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4466 & _GEN_3977) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_31_line_3 <= _GEN_2946;
        end else begin
          cache_31_line_3 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_31_line_3 <= _GEN_2143;
      end
    end else begin
      cache_31_line_3 <= _GEN_2143;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_31_line_4 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4466 & _GEN_3979) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_31_line_4 <= _GEN_2946;
        end else begin
          cache_31_line_4 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_31_line_4 <= _GEN_2207;
      end
    end else begin
      cache_31_line_4 <= _GEN_2207;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_31_line_5 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4466 & _GEN_3981) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_31_line_5 <= _GEN_2946;
        end else begin
          cache_31_line_5 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_31_line_5 <= _GEN_2271;
      end
    end else begin
      cache_31_line_5 <= _GEN_2271;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_31_line_6 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4466 & _GEN_3983) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_31_line_6 <= _GEN_2946;
        end else begin
          cache_31_line_6 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_31_line_6 <= _GEN_2335;
      end
    end else begin
      cache_31_line_6 <= _GEN_2335;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_31_line_7 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4466 & _GEN_3985) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_31_line_7 <= _GEN_2946;
        end else begin
          cache_31_line_7 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_31_line_7 <= _GEN_2399;
      end
    end else begin
      cache_31_line_7 <= _GEN_2399;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_32_validBit <= 1'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      cache_32_validBit <= _GEN_1184;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_32_tag <= 5'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      if (6'h20 == cacheLine) begin // @[Cache.scala 50:26]
        cache_32_tag <= tag; // @[Cache.scala 50:26]
      end
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_32_line_0 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4482 & _GEN_3987) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_32_line_0 <= _GEN_2946;
        end else begin
          cache_32_line_0 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_32_line_0 <= _GEN_1952;
      end
    end else begin
      cache_32_line_0 <= _GEN_1952;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_32_line_1 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4482 & _GEN_3973) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_32_line_1 <= _GEN_2946;
        end else begin
          cache_32_line_1 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_32_line_1 <= _GEN_2016;
      end
    end else begin
      cache_32_line_1 <= _GEN_2016;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_32_line_2 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4482 & _GEN_3975) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_32_line_2 <= _GEN_2946;
        end else begin
          cache_32_line_2 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_32_line_2 <= _GEN_2080;
      end
    end else begin
      cache_32_line_2 <= _GEN_2080;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_32_line_3 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4482 & _GEN_3977) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_32_line_3 <= _GEN_2946;
        end else begin
          cache_32_line_3 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_32_line_3 <= _GEN_2144;
      end
    end else begin
      cache_32_line_3 <= _GEN_2144;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_32_line_4 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4482 & _GEN_3979) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_32_line_4 <= _GEN_2946;
        end else begin
          cache_32_line_4 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_32_line_4 <= _GEN_2208;
      end
    end else begin
      cache_32_line_4 <= _GEN_2208;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_32_line_5 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4482 & _GEN_3981) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_32_line_5 <= _GEN_2946;
        end else begin
          cache_32_line_5 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_32_line_5 <= _GEN_2272;
      end
    end else begin
      cache_32_line_5 <= _GEN_2272;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_32_line_6 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4482 & _GEN_3983) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_32_line_6 <= _GEN_2946;
        end else begin
          cache_32_line_6 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_32_line_6 <= _GEN_2336;
      end
    end else begin
      cache_32_line_6 <= _GEN_2336;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_32_line_7 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4482 & _GEN_3985) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_32_line_7 <= _GEN_2946;
        end else begin
          cache_32_line_7 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_32_line_7 <= _GEN_2400;
      end
    end else begin
      cache_32_line_7 <= _GEN_2400;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_33_validBit <= 1'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      cache_33_validBit <= _GEN_1185;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_33_tag <= 5'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      if (6'h21 == cacheLine) begin // @[Cache.scala 50:26]
        cache_33_tag <= tag; // @[Cache.scala 50:26]
      end
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_33_line_0 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4498 & _GEN_3987) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_33_line_0 <= _GEN_2946;
        end else begin
          cache_33_line_0 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_33_line_0 <= _GEN_1953;
      end
    end else begin
      cache_33_line_0 <= _GEN_1953;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_33_line_1 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4498 & _GEN_3973) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_33_line_1 <= _GEN_2946;
        end else begin
          cache_33_line_1 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_33_line_1 <= _GEN_2017;
      end
    end else begin
      cache_33_line_1 <= _GEN_2017;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_33_line_2 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4498 & _GEN_3975) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_33_line_2 <= _GEN_2946;
        end else begin
          cache_33_line_2 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_33_line_2 <= _GEN_2081;
      end
    end else begin
      cache_33_line_2 <= _GEN_2081;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_33_line_3 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4498 & _GEN_3977) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_33_line_3 <= _GEN_2946;
        end else begin
          cache_33_line_3 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_33_line_3 <= _GEN_2145;
      end
    end else begin
      cache_33_line_3 <= _GEN_2145;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_33_line_4 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4498 & _GEN_3979) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_33_line_4 <= _GEN_2946;
        end else begin
          cache_33_line_4 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_33_line_4 <= _GEN_2209;
      end
    end else begin
      cache_33_line_4 <= _GEN_2209;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_33_line_5 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4498 & _GEN_3981) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_33_line_5 <= _GEN_2946;
        end else begin
          cache_33_line_5 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_33_line_5 <= _GEN_2273;
      end
    end else begin
      cache_33_line_5 <= _GEN_2273;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_33_line_6 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4498 & _GEN_3983) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_33_line_6 <= _GEN_2946;
        end else begin
          cache_33_line_6 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_33_line_6 <= _GEN_2337;
      end
    end else begin
      cache_33_line_6 <= _GEN_2337;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_33_line_7 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4498 & _GEN_3985) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_33_line_7 <= _GEN_2946;
        end else begin
          cache_33_line_7 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_33_line_7 <= _GEN_2401;
      end
    end else begin
      cache_33_line_7 <= _GEN_2401;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_34_validBit <= 1'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      cache_34_validBit <= _GEN_1186;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_34_tag <= 5'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      if (6'h22 == cacheLine) begin // @[Cache.scala 50:26]
        cache_34_tag <= tag; // @[Cache.scala 50:26]
      end
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_34_line_0 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4514 & _GEN_3987) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_34_line_0 <= _GEN_2946;
        end else begin
          cache_34_line_0 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_34_line_0 <= _GEN_1954;
      end
    end else begin
      cache_34_line_0 <= _GEN_1954;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_34_line_1 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4514 & _GEN_3973) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_34_line_1 <= _GEN_2946;
        end else begin
          cache_34_line_1 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_34_line_1 <= _GEN_2018;
      end
    end else begin
      cache_34_line_1 <= _GEN_2018;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_34_line_2 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4514 & _GEN_3975) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_34_line_2 <= _GEN_2946;
        end else begin
          cache_34_line_2 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_34_line_2 <= _GEN_2082;
      end
    end else begin
      cache_34_line_2 <= _GEN_2082;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_34_line_3 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4514 & _GEN_3977) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_34_line_3 <= _GEN_2946;
        end else begin
          cache_34_line_3 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_34_line_3 <= _GEN_2146;
      end
    end else begin
      cache_34_line_3 <= _GEN_2146;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_34_line_4 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4514 & _GEN_3979) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_34_line_4 <= _GEN_2946;
        end else begin
          cache_34_line_4 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_34_line_4 <= _GEN_2210;
      end
    end else begin
      cache_34_line_4 <= _GEN_2210;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_34_line_5 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4514 & _GEN_3981) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_34_line_5 <= _GEN_2946;
        end else begin
          cache_34_line_5 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_34_line_5 <= _GEN_2274;
      end
    end else begin
      cache_34_line_5 <= _GEN_2274;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_34_line_6 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4514 & _GEN_3983) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_34_line_6 <= _GEN_2946;
        end else begin
          cache_34_line_6 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_34_line_6 <= _GEN_2338;
      end
    end else begin
      cache_34_line_6 <= _GEN_2338;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_34_line_7 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4514 & _GEN_3985) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_34_line_7 <= _GEN_2946;
        end else begin
          cache_34_line_7 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_34_line_7 <= _GEN_2402;
      end
    end else begin
      cache_34_line_7 <= _GEN_2402;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_35_validBit <= 1'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      cache_35_validBit <= _GEN_1187;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_35_tag <= 5'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      if (6'h23 == cacheLine) begin // @[Cache.scala 50:26]
        cache_35_tag <= tag; // @[Cache.scala 50:26]
      end
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_35_line_0 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4530 & _GEN_3987) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_35_line_0 <= _GEN_2946;
        end else begin
          cache_35_line_0 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_35_line_0 <= _GEN_1955;
      end
    end else begin
      cache_35_line_0 <= _GEN_1955;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_35_line_1 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4530 & _GEN_3973) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_35_line_1 <= _GEN_2946;
        end else begin
          cache_35_line_1 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_35_line_1 <= _GEN_2019;
      end
    end else begin
      cache_35_line_1 <= _GEN_2019;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_35_line_2 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4530 & _GEN_3975) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_35_line_2 <= _GEN_2946;
        end else begin
          cache_35_line_2 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_35_line_2 <= _GEN_2083;
      end
    end else begin
      cache_35_line_2 <= _GEN_2083;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_35_line_3 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4530 & _GEN_3977) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_35_line_3 <= _GEN_2946;
        end else begin
          cache_35_line_3 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_35_line_3 <= _GEN_2147;
      end
    end else begin
      cache_35_line_3 <= _GEN_2147;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_35_line_4 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4530 & _GEN_3979) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_35_line_4 <= _GEN_2946;
        end else begin
          cache_35_line_4 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_35_line_4 <= _GEN_2211;
      end
    end else begin
      cache_35_line_4 <= _GEN_2211;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_35_line_5 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4530 & _GEN_3981) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_35_line_5 <= _GEN_2946;
        end else begin
          cache_35_line_5 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_35_line_5 <= _GEN_2275;
      end
    end else begin
      cache_35_line_5 <= _GEN_2275;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_35_line_6 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4530 & _GEN_3983) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_35_line_6 <= _GEN_2946;
        end else begin
          cache_35_line_6 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_35_line_6 <= _GEN_2339;
      end
    end else begin
      cache_35_line_6 <= _GEN_2339;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_35_line_7 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4530 & _GEN_3985) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_35_line_7 <= _GEN_2946;
        end else begin
          cache_35_line_7 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_35_line_7 <= _GEN_2403;
      end
    end else begin
      cache_35_line_7 <= _GEN_2403;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_36_validBit <= 1'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      cache_36_validBit <= _GEN_1188;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_36_tag <= 5'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      if (6'h24 == cacheLine) begin // @[Cache.scala 50:26]
        cache_36_tag <= tag; // @[Cache.scala 50:26]
      end
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_36_line_0 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4546 & _GEN_3987) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_36_line_0 <= _GEN_2946;
        end else begin
          cache_36_line_0 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_36_line_0 <= _GEN_1956;
      end
    end else begin
      cache_36_line_0 <= _GEN_1956;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_36_line_1 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4546 & _GEN_3973) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_36_line_1 <= _GEN_2946;
        end else begin
          cache_36_line_1 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_36_line_1 <= _GEN_2020;
      end
    end else begin
      cache_36_line_1 <= _GEN_2020;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_36_line_2 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4546 & _GEN_3975) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_36_line_2 <= _GEN_2946;
        end else begin
          cache_36_line_2 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_36_line_2 <= _GEN_2084;
      end
    end else begin
      cache_36_line_2 <= _GEN_2084;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_36_line_3 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4546 & _GEN_3977) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_36_line_3 <= _GEN_2946;
        end else begin
          cache_36_line_3 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_36_line_3 <= _GEN_2148;
      end
    end else begin
      cache_36_line_3 <= _GEN_2148;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_36_line_4 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4546 & _GEN_3979) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_36_line_4 <= _GEN_2946;
        end else begin
          cache_36_line_4 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_36_line_4 <= _GEN_2212;
      end
    end else begin
      cache_36_line_4 <= _GEN_2212;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_36_line_5 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4546 & _GEN_3981) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_36_line_5 <= _GEN_2946;
        end else begin
          cache_36_line_5 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_36_line_5 <= _GEN_2276;
      end
    end else begin
      cache_36_line_5 <= _GEN_2276;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_36_line_6 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4546 & _GEN_3983) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_36_line_6 <= _GEN_2946;
        end else begin
          cache_36_line_6 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_36_line_6 <= _GEN_2340;
      end
    end else begin
      cache_36_line_6 <= _GEN_2340;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_36_line_7 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4546 & _GEN_3985) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_36_line_7 <= _GEN_2946;
        end else begin
          cache_36_line_7 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_36_line_7 <= _GEN_2404;
      end
    end else begin
      cache_36_line_7 <= _GEN_2404;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_37_validBit <= 1'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      cache_37_validBit <= _GEN_1189;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_37_tag <= 5'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      if (6'h25 == cacheLine) begin // @[Cache.scala 50:26]
        cache_37_tag <= tag; // @[Cache.scala 50:26]
      end
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_37_line_0 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4562 & _GEN_3987) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_37_line_0 <= _GEN_2946;
        end else begin
          cache_37_line_0 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_37_line_0 <= _GEN_1957;
      end
    end else begin
      cache_37_line_0 <= _GEN_1957;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_37_line_1 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4562 & _GEN_3973) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_37_line_1 <= _GEN_2946;
        end else begin
          cache_37_line_1 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_37_line_1 <= _GEN_2021;
      end
    end else begin
      cache_37_line_1 <= _GEN_2021;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_37_line_2 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4562 & _GEN_3975) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_37_line_2 <= _GEN_2946;
        end else begin
          cache_37_line_2 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_37_line_2 <= _GEN_2085;
      end
    end else begin
      cache_37_line_2 <= _GEN_2085;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_37_line_3 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4562 & _GEN_3977) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_37_line_3 <= _GEN_2946;
        end else begin
          cache_37_line_3 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_37_line_3 <= _GEN_2149;
      end
    end else begin
      cache_37_line_3 <= _GEN_2149;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_37_line_4 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4562 & _GEN_3979) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_37_line_4 <= _GEN_2946;
        end else begin
          cache_37_line_4 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_37_line_4 <= _GEN_2213;
      end
    end else begin
      cache_37_line_4 <= _GEN_2213;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_37_line_5 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4562 & _GEN_3981) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_37_line_5 <= _GEN_2946;
        end else begin
          cache_37_line_5 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_37_line_5 <= _GEN_2277;
      end
    end else begin
      cache_37_line_5 <= _GEN_2277;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_37_line_6 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4562 & _GEN_3983) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_37_line_6 <= _GEN_2946;
        end else begin
          cache_37_line_6 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_37_line_6 <= _GEN_2341;
      end
    end else begin
      cache_37_line_6 <= _GEN_2341;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_37_line_7 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4562 & _GEN_3985) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_37_line_7 <= _GEN_2946;
        end else begin
          cache_37_line_7 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_37_line_7 <= _GEN_2405;
      end
    end else begin
      cache_37_line_7 <= _GEN_2405;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_38_validBit <= 1'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      cache_38_validBit <= _GEN_1190;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_38_tag <= 5'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      if (6'h26 == cacheLine) begin // @[Cache.scala 50:26]
        cache_38_tag <= tag; // @[Cache.scala 50:26]
      end
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_38_line_0 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4578 & _GEN_3987) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_38_line_0 <= _GEN_2946;
        end else begin
          cache_38_line_0 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_38_line_0 <= _GEN_1958;
      end
    end else begin
      cache_38_line_0 <= _GEN_1958;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_38_line_1 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4578 & _GEN_3973) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_38_line_1 <= _GEN_2946;
        end else begin
          cache_38_line_1 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_38_line_1 <= _GEN_2022;
      end
    end else begin
      cache_38_line_1 <= _GEN_2022;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_38_line_2 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4578 & _GEN_3975) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_38_line_2 <= _GEN_2946;
        end else begin
          cache_38_line_2 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_38_line_2 <= _GEN_2086;
      end
    end else begin
      cache_38_line_2 <= _GEN_2086;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_38_line_3 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4578 & _GEN_3977) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_38_line_3 <= _GEN_2946;
        end else begin
          cache_38_line_3 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_38_line_3 <= _GEN_2150;
      end
    end else begin
      cache_38_line_3 <= _GEN_2150;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_38_line_4 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4578 & _GEN_3979) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_38_line_4 <= _GEN_2946;
        end else begin
          cache_38_line_4 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_38_line_4 <= _GEN_2214;
      end
    end else begin
      cache_38_line_4 <= _GEN_2214;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_38_line_5 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4578 & _GEN_3981) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_38_line_5 <= _GEN_2946;
        end else begin
          cache_38_line_5 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_38_line_5 <= _GEN_2278;
      end
    end else begin
      cache_38_line_5 <= _GEN_2278;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_38_line_6 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4578 & _GEN_3983) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_38_line_6 <= _GEN_2946;
        end else begin
          cache_38_line_6 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_38_line_6 <= _GEN_2342;
      end
    end else begin
      cache_38_line_6 <= _GEN_2342;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_38_line_7 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4578 & _GEN_3985) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_38_line_7 <= _GEN_2946;
        end else begin
          cache_38_line_7 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_38_line_7 <= _GEN_2406;
      end
    end else begin
      cache_38_line_7 <= _GEN_2406;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_39_validBit <= 1'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      cache_39_validBit <= _GEN_1191;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_39_tag <= 5'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      if (6'h27 == cacheLine) begin // @[Cache.scala 50:26]
        cache_39_tag <= tag; // @[Cache.scala 50:26]
      end
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_39_line_0 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4594 & _GEN_3987) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_39_line_0 <= _GEN_2946;
        end else begin
          cache_39_line_0 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_39_line_0 <= _GEN_1959;
      end
    end else begin
      cache_39_line_0 <= _GEN_1959;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_39_line_1 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4594 & _GEN_3973) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_39_line_1 <= _GEN_2946;
        end else begin
          cache_39_line_1 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_39_line_1 <= _GEN_2023;
      end
    end else begin
      cache_39_line_1 <= _GEN_2023;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_39_line_2 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4594 & _GEN_3975) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_39_line_2 <= _GEN_2946;
        end else begin
          cache_39_line_2 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_39_line_2 <= _GEN_2087;
      end
    end else begin
      cache_39_line_2 <= _GEN_2087;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_39_line_3 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4594 & _GEN_3977) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_39_line_3 <= _GEN_2946;
        end else begin
          cache_39_line_3 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_39_line_3 <= _GEN_2151;
      end
    end else begin
      cache_39_line_3 <= _GEN_2151;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_39_line_4 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4594 & _GEN_3979) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_39_line_4 <= _GEN_2946;
        end else begin
          cache_39_line_4 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_39_line_4 <= _GEN_2215;
      end
    end else begin
      cache_39_line_4 <= _GEN_2215;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_39_line_5 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4594 & _GEN_3981) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_39_line_5 <= _GEN_2946;
        end else begin
          cache_39_line_5 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_39_line_5 <= _GEN_2279;
      end
    end else begin
      cache_39_line_5 <= _GEN_2279;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_39_line_6 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4594 & _GEN_3983) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_39_line_6 <= _GEN_2946;
        end else begin
          cache_39_line_6 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_39_line_6 <= _GEN_2343;
      end
    end else begin
      cache_39_line_6 <= _GEN_2343;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_39_line_7 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4594 & _GEN_3985) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_39_line_7 <= _GEN_2946;
        end else begin
          cache_39_line_7 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_39_line_7 <= _GEN_2407;
      end
    end else begin
      cache_39_line_7 <= _GEN_2407;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_40_validBit <= 1'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      cache_40_validBit <= _GEN_1192;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_40_tag <= 5'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      if (6'h28 == cacheLine) begin // @[Cache.scala 50:26]
        cache_40_tag <= tag; // @[Cache.scala 50:26]
      end
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_40_line_0 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4610 & _GEN_3987) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_40_line_0 <= _GEN_2946;
        end else begin
          cache_40_line_0 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_40_line_0 <= _GEN_1960;
      end
    end else begin
      cache_40_line_0 <= _GEN_1960;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_40_line_1 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4610 & _GEN_3973) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_40_line_1 <= _GEN_2946;
        end else begin
          cache_40_line_1 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_40_line_1 <= _GEN_2024;
      end
    end else begin
      cache_40_line_1 <= _GEN_2024;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_40_line_2 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4610 & _GEN_3975) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_40_line_2 <= _GEN_2946;
        end else begin
          cache_40_line_2 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_40_line_2 <= _GEN_2088;
      end
    end else begin
      cache_40_line_2 <= _GEN_2088;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_40_line_3 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4610 & _GEN_3977) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_40_line_3 <= _GEN_2946;
        end else begin
          cache_40_line_3 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_40_line_3 <= _GEN_2152;
      end
    end else begin
      cache_40_line_3 <= _GEN_2152;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_40_line_4 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4610 & _GEN_3979) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_40_line_4 <= _GEN_2946;
        end else begin
          cache_40_line_4 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_40_line_4 <= _GEN_2216;
      end
    end else begin
      cache_40_line_4 <= _GEN_2216;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_40_line_5 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4610 & _GEN_3981) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_40_line_5 <= _GEN_2946;
        end else begin
          cache_40_line_5 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_40_line_5 <= _GEN_2280;
      end
    end else begin
      cache_40_line_5 <= _GEN_2280;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_40_line_6 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4610 & _GEN_3983) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_40_line_6 <= _GEN_2946;
        end else begin
          cache_40_line_6 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_40_line_6 <= _GEN_2344;
      end
    end else begin
      cache_40_line_6 <= _GEN_2344;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_40_line_7 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4610 & _GEN_3985) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_40_line_7 <= _GEN_2946;
        end else begin
          cache_40_line_7 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_40_line_7 <= _GEN_2408;
      end
    end else begin
      cache_40_line_7 <= _GEN_2408;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_41_validBit <= 1'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      cache_41_validBit <= _GEN_1193;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_41_tag <= 5'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      if (6'h29 == cacheLine) begin // @[Cache.scala 50:26]
        cache_41_tag <= tag; // @[Cache.scala 50:26]
      end
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_41_line_0 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4626 & _GEN_3987) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_41_line_0 <= _GEN_2946;
        end else begin
          cache_41_line_0 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_41_line_0 <= _GEN_1961;
      end
    end else begin
      cache_41_line_0 <= _GEN_1961;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_41_line_1 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4626 & _GEN_3973) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_41_line_1 <= _GEN_2946;
        end else begin
          cache_41_line_1 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_41_line_1 <= _GEN_2025;
      end
    end else begin
      cache_41_line_1 <= _GEN_2025;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_41_line_2 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4626 & _GEN_3975) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_41_line_2 <= _GEN_2946;
        end else begin
          cache_41_line_2 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_41_line_2 <= _GEN_2089;
      end
    end else begin
      cache_41_line_2 <= _GEN_2089;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_41_line_3 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4626 & _GEN_3977) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_41_line_3 <= _GEN_2946;
        end else begin
          cache_41_line_3 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_41_line_3 <= _GEN_2153;
      end
    end else begin
      cache_41_line_3 <= _GEN_2153;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_41_line_4 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4626 & _GEN_3979) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_41_line_4 <= _GEN_2946;
        end else begin
          cache_41_line_4 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_41_line_4 <= _GEN_2217;
      end
    end else begin
      cache_41_line_4 <= _GEN_2217;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_41_line_5 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4626 & _GEN_3981) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_41_line_5 <= _GEN_2946;
        end else begin
          cache_41_line_5 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_41_line_5 <= _GEN_2281;
      end
    end else begin
      cache_41_line_5 <= _GEN_2281;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_41_line_6 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4626 & _GEN_3983) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_41_line_6 <= _GEN_2946;
        end else begin
          cache_41_line_6 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_41_line_6 <= _GEN_2345;
      end
    end else begin
      cache_41_line_6 <= _GEN_2345;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_41_line_7 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4626 & _GEN_3985) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_41_line_7 <= _GEN_2946;
        end else begin
          cache_41_line_7 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_41_line_7 <= _GEN_2409;
      end
    end else begin
      cache_41_line_7 <= _GEN_2409;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_42_validBit <= 1'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      cache_42_validBit <= _GEN_1194;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_42_tag <= 5'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      if (6'h2a == cacheLine) begin // @[Cache.scala 50:26]
        cache_42_tag <= tag; // @[Cache.scala 50:26]
      end
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_42_line_0 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4642 & _GEN_3987) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_42_line_0 <= _GEN_2946;
        end else begin
          cache_42_line_0 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_42_line_0 <= _GEN_1962;
      end
    end else begin
      cache_42_line_0 <= _GEN_1962;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_42_line_1 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4642 & _GEN_3973) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_42_line_1 <= _GEN_2946;
        end else begin
          cache_42_line_1 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_42_line_1 <= _GEN_2026;
      end
    end else begin
      cache_42_line_1 <= _GEN_2026;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_42_line_2 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4642 & _GEN_3975) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_42_line_2 <= _GEN_2946;
        end else begin
          cache_42_line_2 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_42_line_2 <= _GEN_2090;
      end
    end else begin
      cache_42_line_2 <= _GEN_2090;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_42_line_3 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4642 & _GEN_3977) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_42_line_3 <= _GEN_2946;
        end else begin
          cache_42_line_3 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_42_line_3 <= _GEN_2154;
      end
    end else begin
      cache_42_line_3 <= _GEN_2154;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_42_line_4 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4642 & _GEN_3979) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_42_line_4 <= _GEN_2946;
        end else begin
          cache_42_line_4 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_42_line_4 <= _GEN_2218;
      end
    end else begin
      cache_42_line_4 <= _GEN_2218;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_42_line_5 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4642 & _GEN_3981) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_42_line_5 <= _GEN_2946;
        end else begin
          cache_42_line_5 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_42_line_5 <= _GEN_2282;
      end
    end else begin
      cache_42_line_5 <= _GEN_2282;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_42_line_6 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4642 & _GEN_3983) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_42_line_6 <= _GEN_2946;
        end else begin
          cache_42_line_6 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_42_line_6 <= _GEN_2346;
      end
    end else begin
      cache_42_line_6 <= _GEN_2346;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_42_line_7 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4642 & _GEN_3985) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_42_line_7 <= _GEN_2946;
        end else begin
          cache_42_line_7 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_42_line_7 <= _GEN_2410;
      end
    end else begin
      cache_42_line_7 <= _GEN_2410;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_43_validBit <= 1'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      cache_43_validBit <= _GEN_1195;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_43_tag <= 5'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      if (6'h2b == cacheLine) begin // @[Cache.scala 50:26]
        cache_43_tag <= tag; // @[Cache.scala 50:26]
      end
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_43_line_0 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4658 & _GEN_3987) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_43_line_0 <= _GEN_2946;
        end else begin
          cache_43_line_0 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_43_line_0 <= _GEN_1963;
      end
    end else begin
      cache_43_line_0 <= _GEN_1963;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_43_line_1 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4658 & _GEN_3973) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_43_line_1 <= _GEN_2946;
        end else begin
          cache_43_line_1 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_43_line_1 <= _GEN_2027;
      end
    end else begin
      cache_43_line_1 <= _GEN_2027;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_43_line_2 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4658 & _GEN_3975) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_43_line_2 <= _GEN_2946;
        end else begin
          cache_43_line_2 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_43_line_2 <= _GEN_2091;
      end
    end else begin
      cache_43_line_2 <= _GEN_2091;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_43_line_3 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4658 & _GEN_3977) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_43_line_3 <= _GEN_2946;
        end else begin
          cache_43_line_3 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_43_line_3 <= _GEN_2155;
      end
    end else begin
      cache_43_line_3 <= _GEN_2155;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_43_line_4 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4658 & _GEN_3979) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_43_line_4 <= _GEN_2946;
        end else begin
          cache_43_line_4 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_43_line_4 <= _GEN_2219;
      end
    end else begin
      cache_43_line_4 <= _GEN_2219;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_43_line_5 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4658 & _GEN_3981) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_43_line_5 <= _GEN_2946;
        end else begin
          cache_43_line_5 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_43_line_5 <= _GEN_2283;
      end
    end else begin
      cache_43_line_5 <= _GEN_2283;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_43_line_6 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4658 & _GEN_3983) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_43_line_6 <= _GEN_2946;
        end else begin
          cache_43_line_6 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_43_line_6 <= _GEN_2347;
      end
    end else begin
      cache_43_line_6 <= _GEN_2347;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_43_line_7 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4658 & _GEN_3985) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_43_line_7 <= _GEN_2946;
        end else begin
          cache_43_line_7 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_43_line_7 <= _GEN_2411;
      end
    end else begin
      cache_43_line_7 <= _GEN_2411;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_44_validBit <= 1'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      cache_44_validBit <= _GEN_1196;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_44_tag <= 5'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      if (6'h2c == cacheLine) begin // @[Cache.scala 50:26]
        cache_44_tag <= tag; // @[Cache.scala 50:26]
      end
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_44_line_0 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4674 & _GEN_3987) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_44_line_0 <= _GEN_2946;
        end else begin
          cache_44_line_0 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_44_line_0 <= _GEN_1964;
      end
    end else begin
      cache_44_line_0 <= _GEN_1964;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_44_line_1 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4674 & _GEN_3973) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_44_line_1 <= _GEN_2946;
        end else begin
          cache_44_line_1 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_44_line_1 <= _GEN_2028;
      end
    end else begin
      cache_44_line_1 <= _GEN_2028;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_44_line_2 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4674 & _GEN_3975) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_44_line_2 <= _GEN_2946;
        end else begin
          cache_44_line_2 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_44_line_2 <= _GEN_2092;
      end
    end else begin
      cache_44_line_2 <= _GEN_2092;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_44_line_3 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4674 & _GEN_3977) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_44_line_3 <= _GEN_2946;
        end else begin
          cache_44_line_3 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_44_line_3 <= _GEN_2156;
      end
    end else begin
      cache_44_line_3 <= _GEN_2156;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_44_line_4 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4674 & _GEN_3979) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_44_line_4 <= _GEN_2946;
        end else begin
          cache_44_line_4 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_44_line_4 <= _GEN_2220;
      end
    end else begin
      cache_44_line_4 <= _GEN_2220;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_44_line_5 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4674 & _GEN_3981) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_44_line_5 <= _GEN_2946;
        end else begin
          cache_44_line_5 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_44_line_5 <= _GEN_2284;
      end
    end else begin
      cache_44_line_5 <= _GEN_2284;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_44_line_6 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4674 & _GEN_3983) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_44_line_6 <= _GEN_2946;
        end else begin
          cache_44_line_6 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_44_line_6 <= _GEN_2348;
      end
    end else begin
      cache_44_line_6 <= _GEN_2348;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_44_line_7 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4674 & _GEN_3985) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_44_line_7 <= _GEN_2946;
        end else begin
          cache_44_line_7 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_44_line_7 <= _GEN_2412;
      end
    end else begin
      cache_44_line_7 <= _GEN_2412;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_45_validBit <= 1'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      cache_45_validBit <= _GEN_1197;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_45_tag <= 5'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      if (6'h2d == cacheLine) begin // @[Cache.scala 50:26]
        cache_45_tag <= tag; // @[Cache.scala 50:26]
      end
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_45_line_0 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4690 & _GEN_3987) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_45_line_0 <= _GEN_2946;
        end else begin
          cache_45_line_0 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_45_line_0 <= _GEN_1965;
      end
    end else begin
      cache_45_line_0 <= _GEN_1965;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_45_line_1 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4690 & _GEN_3973) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_45_line_1 <= _GEN_2946;
        end else begin
          cache_45_line_1 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_45_line_1 <= _GEN_2029;
      end
    end else begin
      cache_45_line_1 <= _GEN_2029;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_45_line_2 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4690 & _GEN_3975) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_45_line_2 <= _GEN_2946;
        end else begin
          cache_45_line_2 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_45_line_2 <= _GEN_2093;
      end
    end else begin
      cache_45_line_2 <= _GEN_2093;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_45_line_3 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4690 & _GEN_3977) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_45_line_3 <= _GEN_2946;
        end else begin
          cache_45_line_3 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_45_line_3 <= _GEN_2157;
      end
    end else begin
      cache_45_line_3 <= _GEN_2157;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_45_line_4 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4690 & _GEN_3979) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_45_line_4 <= _GEN_2946;
        end else begin
          cache_45_line_4 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_45_line_4 <= _GEN_2221;
      end
    end else begin
      cache_45_line_4 <= _GEN_2221;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_45_line_5 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4690 & _GEN_3981) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_45_line_5 <= _GEN_2946;
        end else begin
          cache_45_line_5 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_45_line_5 <= _GEN_2285;
      end
    end else begin
      cache_45_line_5 <= _GEN_2285;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_45_line_6 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4690 & _GEN_3983) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_45_line_6 <= _GEN_2946;
        end else begin
          cache_45_line_6 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_45_line_6 <= _GEN_2349;
      end
    end else begin
      cache_45_line_6 <= _GEN_2349;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_45_line_7 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4690 & _GEN_3985) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_45_line_7 <= _GEN_2946;
        end else begin
          cache_45_line_7 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_45_line_7 <= _GEN_2413;
      end
    end else begin
      cache_45_line_7 <= _GEN_2413;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_46_validBit <= 1'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      cache_46_validBit <= _GEN_1198;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_46_tag <= 5'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      if (6'h2e == cacheLine) begin // @[Cache.scala 50:26]
        cache_46_tag <= tag; // @[Cache.scala 50:26]
      end
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_46_line_0 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4706 & _GEN_3987) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_46_line_0 <= _GEN_2946;
        end else begin
          cache_46_line_0 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_46_line_0 <= _GEN_1966;
      end
    end else begin
      cache_46_line_0 <= _GEN_1966;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_46_line_1 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4706 & _GEN_3973) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_46_line_1 <= _GEN_2946;
        end else begin
          cache_46_line_1 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_46_line_1 <= _GEN_2030;
      end
    end else begin
      cache_46_line_1 <= _GEN_2030;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_46_line_2 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4706 & _GEN_3975) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_46_line_2 <= _GEN_2946;
        end else begin
          cache_46_line_2 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_46_line_2 <= _GEN_2094;
      end
    end else begin
      cache_46_line_2 <= _GEN_2094;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_46_line_3 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4706 & _GEN_3977) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_46_line_3 <= _GEN_2946;
        end else begin
          cache_46_line_3 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_46_line_3 <= _GEN_2158;
      end
    end else begin
      cache_46_line_3 <= _GEN_2158;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_46_line_4 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4706 & _GEN_3979) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_46_line_4 <= _GEN_2946;
        end else begin
          cache_46_line_4 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_46_line_4 <= _GEN_2222;
      end
    end else begin
      cache_46_line_4 <= _GEN_2222;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_46_line_5 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4706 & _GEN_3981) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_46_line_5 <= _GEN_2946;
        end else begin
          cache_46_line_5 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_46_line_5 <= _GEN_2286;
      end
    end else begin
      cache_46_line_5 <= _GEN_2286;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_46_line_6 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4706 & _GEN_3983) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_46_line_6 <= _GEN_2946;
        end else begin
          cache_46_line_6 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_46_line_6 <= _GEN_2350;
      end
    end else begin
      cache_46_line_6 <= _GEN_2350;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_46_line_7 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4706 & _GEN_3985) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_46_line_7 <= _GEN_2946;
        end else begin
          cache_46_line_7 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_46_line_7 <= _GEN_2414;
      end
    end else begin
      cache_46_line_7 <= _GEN_2414;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_47_validBit <= 1'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      cache_47_validBit <= _GEN_1199;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_47_tag <= 5'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      if (6'h2f == cacheLine) begin // @[Cache.scala 50:26]
        cache_47_tag <= tag; // @[Cache.scala 50:26]
      end
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_47_line_0 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4722 & _GEN_3987) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_47_line_0 <= _GEN_2946;
        end else begin
          cache_47_line_0 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_47_line_0 <= _GEN_1967;
      end
    end else begin
      cache_47_line_0 <= _GEN_1967;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_47_line_1 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4722 & _GEN_3973) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_47_line_1 <= _GEN_2946;
        end else begin
          cache_47_line_1 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_47_line_1 <= _GEN_2031;
      end
    end else begin
      cache_47_line_1 <= _GEN_2031;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_47_line_2 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4722 & _GEN_3975) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_47_line_2 <= _GEN_2946;
        end else begin
          cache_47_line_2 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_47_line_2 <= _GEN_2095;
      end
    end else begin
      cache_47_line_2 <= _GEN_2095;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_47_line_3 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4722 & _GEN_3977) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_47_line_3 <= _GEN_2946;
        end else begin
          cache_47_line_3 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_47_line_3 <= _GEN_2159;
      end
    end else begin
      cache_47_line_3 <= _GEN_2159;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_47_line_4 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4722 & _GEN_3979) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_47_line_4 <= _GEN_2946;
        end else begin
          cache_47_line_4 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_47_line_4 <= _GEN_2223;
      end
    end else begin
      cache_47_line_4 <= _GEN_2223;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_47_line_5 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4722 & _GEN_3981) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_47_line_5 <= _GEN_2946;
        end else begin
          cache_47_line_5 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_47_line_5 <= _GEN_2287;
      end
    end else begin
      cache_47_line_5 <= _GEN_2287;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_47_line_6 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4722 & _GEN_3983) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_47_line_6 <= _GEN_2946;
        end else begin
          cache_47_line_6 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_47_line_6 <= _GEN_2351;
      end
    end else begin
      cache_47_line_6 <= _GEN_2351;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_47_line_7 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4722 & _GEN_3985) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_47_line_7 <= _GEN_2946;
        end else begin
          cache_47_line_7 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_47_line_7 <= _GEN_2415;
      end
    end else begin
      cache_47_line_7 <= _GEN_2415;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_48_validBit <= 1'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      cache_48_validBit <= _GEN_1200;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_48_tag <= 5'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      if (6'h30 == cacheLine) begin // @[Cache.scala 50:26]
        cache_48_tag <= tag; // @[Cache.scala 50:26]
      end
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_48_line_0 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4738 & _GEN_3987) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_48_line_0 <= _GEN_2946;
        end else begin
          cache_48_line_0 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_48_line_0 <= _GEN_1968;
      end
    end else begin
      cache_48_line_0 <= _GEN_1968;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_48_line_1 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4738 & _GEN_3973) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_48_line_1 <= _GEN_2946;
        end else begin
          cache_48_line_1 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_48_line_1 <= _GEN_2032;
      end
    end else begin
      cache_48_line_1 <= _GEN_2032;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_48_line_2 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4738 & _GEN_3975) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_48_line_2 <= _GEN_2946;
        end else begin
          cache_48_line_2 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_48_line_2 <= _GEN_2096;
      end
    end else begin
      cache_48_line_2 <= _GEN_2096;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_48_line_3 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4738 & _GEN_3977) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_48_line_3 <= _GEN_2946;
        end else begin
          cache_48_line_3 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_48_line_3 <= _GEN_2160;
      end
    end else begin
      cache_48_line_3 <= _GEN_2160;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_48_line_4 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4738 & _GEN_3979) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_48_line_4 <= _GEN_2946;
        end else begin
          cache_48_line_4 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_48_line_4 <= _GEN_2224;
      end
    end else begin
      cache_48_line_4 <= _GEN_2224;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_48_line_5 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4738 & _GEN_3981) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_48_line_5 <= _GEN_2946;
        end else begin
          cache_48_line_5 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_48_line_5 <= _GEN_2288;
      end
    end else begin
      cache_48_line_5 <= _GEN_2288;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_48_line_6 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4738 & _GEN_3983) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_48_line_6 <= _GEN_2946;
        end else begin
          cache_48_line_6 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_48_line_6 <= _GEN_2352;
      end
    end else begin
      cache_48_line_6 <= _GEN_2352;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_48_line_7 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4738 & _GEN_3985) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_48_line_7 <= _GEN_2946;
        end else begin
          cache_48_line_7 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_48_line_7 <= _GEN_2416;
      end
    end else begin
      cache_48_line_7 <= _GEN_2416;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_49_validBit <= 1'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      cache_49_validBit <= _GEN_1201;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_49_tag <= 5'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      if (6'h31 == cacheLine) begin // @[Cache.scala 50:26]
        cache_49_tag <= tag; // @[Cache.scala 50:26]
      end
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_49_line_0 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4754 & _GEN_3987) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_49_line_0 <= _GEN_2946;
        end else begin
          cache_49_line_0 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_49_line_0 <= _GEN_1969;
      end
    end else begin
      cache_49_line_0 <= _GEN_1969;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_49_line_1 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4754 & _GEN_3973) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_49_line_1 <= _GEN_2946;
        end else begin
          cache_49_line_1 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_49_line_1 <= _GEN_2033;
      end
    end else begin
      cache_49_line_1 <= _GEN_2033;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_49_line_2 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4754 & _GEN_3975) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_49_line_2 <= _GEN_2946;
        end else begin
          cache_49_line_2 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_49_line_2 <= _GEN_2097;
      end
    end else begin
      cache_49_line_2 <= _GEN_2097;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_49_line_3 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4754 & _GEN_3977) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_49_line_3 <= _GEN_2946;
        end else begin
          cache_49_line_3 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_49_line_3 <= _GEN_2161;
      end
    end else begin
      cache_49_line_3 <= _GEN_2161;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_49_line_4 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4754 & _GEN_3979) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_49_line_4 <= _GEN_2946;
        end else begin
          cache_49_line_4 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_49_line_4 <= _GEN_2225;
      end
    end else begin
      cache_49_line_4 <= _GEN_2225;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_49_line_5 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4754 & _GEN_3981) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_49_line_5 <= _GEN_2946;
        end else begin
          cache_49_line_5 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_49_line_5 <= _GEN_2289;
      end
    end else begin
      cache_49_line_5 <= _GEN_2289;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_49_line_6 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4754 & _GEN_3983) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_49_line_6 <= _GEN_2946;
        end else begin
          cache_49_line_6 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_49_line_6 <= _GEN_2353;
      end
    end else begin
      cache_49_line_6 <= _GEN_2353;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_49_line_7 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4754 & _GEN_3985) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_49_line_7 <= _GEN_2946;
        end else begin
          cache_49_line_7 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_49_line_7 <= _GEN_2417;
      end
    end else begin
      cache_49_line_7 <= _GEN_2417;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_50_validBit <= 1'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      cache_50_validBit <= _GEN_1202;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_50_tag <= 5'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      if (6'h32 == cacheLine) begin // @[Cache.scala 50:26]
        cache_50_tag <= tag; // @[Cache.scala 50:26]
      end
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_50_line_0 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4770 & _GEN_3987) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_50_line_0 <= _GEN_2946;
        end else begin
          cache_50_line_0 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_50_line_0 <= _GEN_1970;
      end
    end else begin
      cache_50_line_0 <= _GEN_1970;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_50_line_1 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4770 & _GEN_3973) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_50_line_1 <= _GEN_2946;
        end else begin
          cache_50_line_1 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_50_line_1 <= _GEN_2034;
      end
    end else begin
      cache_50_line_1 <= _GEN_2034;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_50_line_2 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4770 & _GEN_3975) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_50_line_2 <= _GEN_2946;
        end else begin
          cache_50_line_2 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_50_line_2 <= _GEN_2098;
      end
    end else begin
      cache_50_line_2 <= _GEN_2098;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_50_line_3 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4770 & _GEN_3977) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_50_line_3 <= _GEN_2946;
        end else begin
          cache_50_line_3 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_50_line_3 <= _GEN_2162;
      end
    end else begin
      cache_50_line_3 <= _GEN_2162;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_50_line_4 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4770 & _GEN_3979) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_50_line_4 <= _GEN_2946;
        end else begin
          cache_50_line_4 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_50_line_4 <= _GEN_2226;
      end
    end else begin
      cache_50_line_4 <= _GEN_2226;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_50_line_5 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4770 & _GEN_3981) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_50_line_5 <= _GEN_2946;
        end else begin
          cache_50_line_5 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_50_line_5 <= _GEN_2290;
      end
    end else begin
      cache_50_line_5 <= _GEN_2290;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_50_line_6 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4770 & _GEN_3983) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_50_line_6 <= _GEN_2946;
        end else begin
          cache_50_line_6 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_50_line_6 <= _GEN_2354;
      end
    end else begin
      cache_50_line_6 <= _GEN_2354;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_50_line_7 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4770 & _GEN_3985) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_50_line_7 <= _GEN_2946;
        end else begin
          cache_50_line_7 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_50_line_7 <= _GEN_2418;
      end
    end else begin
      cache_50_line_7 <= _GEN_2418;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_51_validBit <= 1'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      cache_51_validBit <= _GEN_1203;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_51_tag <= 5'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      if (6'h33 == cacheLine) begin // @[Cache.scala 50:26]
        cache_51_tag <= tag; // @[Cache.scala 50:26]
      end
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_51_line_0 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4786 & _GEN_3987) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_51_line_0 <= _GEN_2946;
        end else begin
          cache_51_line_0 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_51_line_0 <= _GEN_1971;
      end
    end else begin
      cache_51_line_0 <= _GEN_1971;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_51_line_1 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4786 & _GEN_3973) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_51_line_1 <= _GEN_2946;
        end else begin
          cache_51_line_1 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_51_line_1 <= _GEN_2035;
      end
    end else begin
      cache_51_line_1 <= _GEN_2035;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_51_line_2 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4786 & _GEN_3975) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_51_line_2 <= _GEN_2946;
        end else begin
          cache_51_line_2 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_51_line_2 <= _GEN_2099;
      end
    end else begin
      cache_51_line_2 <= _GEN_2099;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_51_line_3 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4786 & _GEN_3977) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_51_line_3 <= _GEN_2946;
        end else begin
          cache_51_line_3 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_51_line_3 <= _GEN_2163;
      end
    end else begin
      cache_51_line_3 <= _GEN_2163;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_51_line_4 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4786 & _GEN_3979) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_51_line_4 <= _GEN_2946;
        end else begin
          cache_51_line_4 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_51_line_4 <= _GEN_2227;
      end
    end else begin
      cache_51_line_4 <= _GEN_2227;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_51_line_5 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4786 & _GEN_3981) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_51_line_5 <= _GEN_2946;
        end else begin
          cache_51_line_5 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_51_line_5 <= _GEN_2291;
      end
    end else begin
      cache_51_line_5 <= _GEN_2291;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_51_line_6 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4786 & _GEN_3983) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_51_line_6 <= _GEN_2946;
        end else begin
          cache_51_line_6 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_51_line_6 <= _GEN_2355;
      end
    end else begin
      cache_51_line_6 <= _GEN_2355;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_51_line_7 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4786 & _GEN_3985) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_51_line_7 <= _GEN_2946;
        end else begin
          cache_51_line_7 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_51_line_7 <= _GEN_2419;
      end
    end else begin
      cache_51_line_7 <= _GEN_2419;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_52_validBit <= 1'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      cache_52_validBit <= _GEN_1204;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_52_tag <= 5'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      if (6'h34 == cacheLine) begin // @[Cache.scala 50:26]
        cache_52_tag <= tag; // @[Cache.scala 50:26]
      end
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_52_line_0 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4802 & _GEN_3987) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_52_line_0 <= _GEN_2946;
        end else begin
          cache_52_line_0 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_52_line_0 <= _GEN_1972;
      end
    end else begin
      cache_52_line_0 <= _GEN_1972;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_52_line_1 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4802 & _GEN_3973) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_52_line_1 <= _GEN_2946;
        end else begin
          cache_52_line_1 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_52_line_1 <= _GEN_2036;
      end
    end else begin
      cache_52_line_1 <= _GEN_2036;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_52_line_2 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4802 & _GEN_3975) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_52_line_2 <= _GEN_2946;
        end else begin
          cache_52_line_2 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_52_line_2 <= _GEN_2100;
      end
    end else begin
      cache_52_line_2 <= _GEN_2100;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_52_line_3 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4802 & _GEN_3977) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_52_line_3 <= _GEN_2946;
        end else begin
          cache_52_line_3 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_52_line_3 <= _GEN_2164;
      end
    end else begin
      cache_52_line_3 <= _GEN_2164;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_52_line_4 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4802 & _GEN_3979) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_52_line_4 <= _GEN_2946;
        end else begin
          cache_52_line_4 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_52_line_4 <= _GEN_2228;
      end
    end else begin
      cache_52_line_4 <= _GEN_2228;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_52_line_5 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4802 & _GEN_3981) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_52_line_5 <= _GEN_2946;
        end else begin
          cache_52_line_5 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_52_line_5 <= _GEN_2292;
      end
    end else begin
      cache_52_line_5 <= _GEN_2292;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_52_line_6 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4802 & _GEN_3983) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_52_line_6 <= _GEN_2946;
        end else begin
          cache_52_line_6 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_52_line_6 <= _GEN_2356;
      end
    end else begin
      cache_52_line_6 <= _GEN_2356;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_52_line_7 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4802 & _GEN_3985) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_52_line_7 <= _GEN_2946;
        end else begin
          cache_52_line_7 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_52_line_7 <= _GEN_2420;
      end
    end else begin
      cache_52_line_7 <= _GEN_2420;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_53_validBit <= 1'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      cache_53_validBit <= _GEN_1205;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_53_tag <= 5'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      if (6'h35 == cacheLine) begin // @[Cache.scala 50:26]
        cache_53_tag <= tag; // @[Cache.scala 50:26]
      end
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_53_line_0 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4818 & _GEN_3987) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_53_line_0 <= _GEN_2946;
        end else begin
          cache_53_line_0 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_53_line_0 <= _GEN_1973;
      end
    end else begin
      cache_53_line_0 <= _GEN_1973;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_53_line_1 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4818 & _GEN_3973) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_53_line_1 <= _GEN_2946;
        end else begin
          cache_53_line_1 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_53_line_1 <= _GEN_2037;
      end
    end else begin
      cache_53_line_1 <= _GEN_2037;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_53_line_2 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4818 & _GEN_3975) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_53_line_2 <= _GEN_2946;
        end else begin
          cache_53_line_2 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_53_line_2 <= _GEN_2101;
      end
    end else begin
      cache_53_line_2 <= _GEN_2101;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_53_line_3 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4818 & _GEN_3977) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_53_line_3 <= _GEN_2946;
        end else begin
          cache_53_line_3 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_53_line_3 <= _GEN_2165;
      end
    end else begin
      cache_53_line_3 <= _GEN_2165;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_53_line_4 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4818 & _GEN_3979) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_53_line_4 <= _GEN_2946;
        end else begin
          cache_53_line_4 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_53_line_4 <= _GEN_2229;
      end
    end else begin
      cache_53_line_4 <= _GEN_2229;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_53_line_5 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4818 & _GEN_3981) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_53_line_5 <= _GEN_2946;
        end else begin
          cache_53_line_5 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_53_line_5 <= _GEN_2293;
      end
    end else begin
      cache_53_line_5 <= _GEN_2293;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_53_line_6 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4818 & _GEN_3983) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_53_line_6 <= _GEN_2946;
        end else begin
          cache_53_line_6 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_53_line_6 <= _GEN_2357;
      end
    end else begin
      cache_53_line_6 <= _GEN_2357;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_53_line_7 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4818 & _GEN_3985) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_53_line_7 <= _GEN_2946;
        end else begin
          cache_53_line_7 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_53_line_7 <= _GEN_2421;
      end
    end else begin
      cache_53_line_7 <= _GEN_2421;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_54_validBit <= 1'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      cache_54_validBit <= _GEN_1206;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_54_tag <= 5'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      if (6'h36 == cacheLine) begin // @[Cache.scala 50:26]
        cache_54_tag <= tag; // @[Cache.scala 50:26]
      end
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_54_line_0 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4834 & _GEN_3987) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_54_line_0 <= _GEN_2946;
        end else begin
          cache_54_line_0 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_54_line_0 <= _GEN_1974;
      end
    end else begin
      cache_54_line_0 <= _GEN_1974;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_54_line_1 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4834 & _GEN_3973) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_54_line_1 <= _GEN_2946;
        end else begin
          cache_54_line_1 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_54_line_1 <= _GEN_2038;
      end
    end else begin
      cache_54_line_1 <= _GEN_2038;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_54_line_2 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4834 & _GEN_3975) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_54_line_2 <= _GEN_2946;
        end else begin
          cache_54_line_2 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_54_line_2 <= _GEN_2102;
      end
    end else begin
      cache_54_line_2 <= _GEN_2102;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_54_line_3 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4834 & _GEN_3977) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_54_line_3 <= _GEN_2946;
        end else begin
          cache_54_line_3 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_54_line_3 <= _GEN_2166;
      end
    end else begin
      cache_54_line_3 <= _GEN_2166;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_54_line_4 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4834 & _GEN_3979) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_54_line_4 <= _GEN_2946;
        end else begin
          cache_54_line_4 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_54_line_4 <= _GEN_2230;
      end
    end else begin
      cache_54_line_4 <= _GEN_2230;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_54_line_5 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4834 & _GEN_3981) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_54_line_5 <= _GEN_2946;
        end else begin
          cache_54_line_5 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_54_line_5 <= _GEN_2294;
      end
    end else begin
      cache_54_line_5 <= _GEN_2294;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_54_line_6 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4834 & _GEN_3983) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_54_line_6 <= _GEN_2946;
        end else begin
          cache_54_line_6 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_54_line_6 <= _GEN_2358;
      end
    end else begin
      cache_54_line_6 <= _GEN_2358;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_54_line_7 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4834 & _GEN_3985) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_54_line_7 <= _GEN_2946;
        end else begin
          cache_54_line_7 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_54_line_7 <= _GEN_2422;
      end
    end else begin
      cache_54_line_7 <= _GEN_2422;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_55_validBit <= 1'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      cache_55_validBit <= _GEN_1207;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_55_tag <= 5'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      if (6'h37 == cacheLine) begin // @[Cache.scala 50:26]
        cache_55_tag <= tag; // @[Cache.scala 50:26]
      end
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_55_line_0 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4850 & _GEN_3987) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_55_line_0 <= _GEN_2946;
        end else begin
          cache_55_line_0 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_55_line_0 <= _GEN_1975;
      end
    end else begin
      cache_55_line_0 <= _GEN_1975;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_55_line_1 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4850 & _GEN_3973) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_55_line_1 <= _GEN_2946;
        end else begin
          cache_55_line_1 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_55_line_1 <= _GEN_2039;
      end
    end else begin
      cache_55_line_1 <= _GEN_2039;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_55_line_2 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4850 & _GEN_3975) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_55_line_2 <= _GEN_2946;
        end else begin
          cache_55_line_2 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_55_line_2 <= _GEN_2103;
      end
    end else begin
      cache_55_line_2 <= _GEN_2103;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_55_line_3 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4850 & _GEN_3977) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_55_line_3 <= _GEN_2946;
        end else begin
          cache_55_line_3 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_55_line_3 <= _GEN_2167;
      end
    end else begin
      cache_55_line_3 <= _GEN_2167;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_55_line_4 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4850 & _GEN_3979) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_55_line_4 <= _GEN_2946;
        end else begin
          cache_55_line_4 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_55_line_4 <= _GEN_2231;
      end
    end else begin
      cache_55_line_4 <= _GEN_2231;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_55_line_5 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4850 & _GEN_3981) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_55_line_5 <= _GEN_2946;
        end else begin
          cache_55_line_5 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_55_line_5 <= _GEN_2295;
      end
    end else begin
      cache_55_line_5 <= _GEN_2295;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_55_line_6 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4850 & _GEN_3983) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_55_line_6 <= _GEN_2946;
        end else begin
          cache_55_line_6 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_55_line_6 <= _GEN_2359;
      end
    end else begin
      cache_55_line_6 <= _GEN_2359;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_55_line_7 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4850 & _GEN_3985) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_55_line_7 <= _GEN_2946;
        end else begin
          cache_55_line_7 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_55_line_7 <= _GEN_2423;
      end
    end else begin
      cache_55_line_7 <= _GEN_2423;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_56_validBit <= 1'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      cache_56_validBit <= _GEN_1208;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_56_tag <= 5'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      if (6'h38 == cacheLine) begin // @[Cache.scala 50:26]
        cache_56_tag <= tag; // @[Cache.scala 50:26]
      end
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_56_line_0 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4866 & _GEN_3987) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_56_line_0 <= _GEN_2946;
        end else begin
          cache_56_line_0 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_56_line_0 <= _GEN_1976;
      end
    end else begin
      cache_56_line_0 <= _GEN_1976;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_56_line_1 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4866 & _GEN_3973) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_56_line_1 <= _GEN_2946;
        end else begin
          cache_56_line_1 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_56_line_1 <= _GEN_2040;
      end
    end else begin
      cache_56_line_1 <= _GEN_2040;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_56_line_2 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4866 & _GEN_3975) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_56_line_2 <= _GEN_2946;
        end else begin
          cache_56_line_2 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_56_line_2 <= _GEN_2104;
      end
    end else begin
      cache_56_line_2 <= _GEN_2104;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_56_line_3 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4866 & _GEN_3977) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_56_line_3 <= _GEN_2946;
        end else begin
          cache_56_line_3 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_56_line_3 <= _GEN_2168;
      end
    end else begin
      cache_56_line_3 <= _GEN_2168;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_56_line_4 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4866 & _GEN_3979) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_56_line_4 <= _GEN_2946;
        end else begin
          cache_56_line_4 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_56_line_4 <= _GEN_2232;
      end
    end else begin
      cache_56_line_4 <= _GEN_2232;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_56_line_5 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4866 & _GEN_3981) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_56_line_5 <= _GEN_2946;
        end else begin
          cache_56_line_5 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_56_line_5 <= _GEN_2296;
      end
    end else begin
      cache_56_line_5 <= _GEN_2296;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_56_line_6 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4866 & _GEN_3983) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_56_line_6 <= _GEN_2946;
        end else begin
          cache_56_line_6 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_56_line_6 <= _GEN_2360;
      end
    end else begin
      cache_56_line_6 <= _GEN_2360;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_56_line_7 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4866 & _GEN_3985) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_56_line_7 <= _GEN_2946;
        end else begin
          cache_56_line_7 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_56_line_7 <= _GEN_2424;
      end
    end else begin
      cache_56_line_7 <= _GEN_2424;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_57_validBit <= 1'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      cache_57_validBit <= _GEN_1209;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_57_tag <= 5'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      if (6'h39 == cacheLine) begin // @[Cache.scala 50:26]
        cache_57_tag <= tag; // @[Cache.scala 50:26]
      end
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_57_line_0 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4882 & _GEN_3987) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_57_line_0 <= _GEN_2946;
        end else begin
          cache_57_line_0 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_57_line_0 <= _GEN_1977;
      end
    end else begin
      cache_57_line_0 <= _GEN_1977;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_57_line_1 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4882 & _GEN_3973) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_57_line_1 <= _GEN_2946;
        end else begin
          cache_57_line_1 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_57_line_1 <= _GEN_2041;
      end
    end else begin
      cache_57_line_1 <= _GEN_2041;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_57_line_2 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4882 & _GEN_3975) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_57_line_2 <= _GEN_2946;
        end else begin
          cache_57_line_2 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_57_line_2 <= _GEN_2105;
      end
    end else begin
      cache_57_line_2 <= _GEN_2105;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_57_line_3 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4882 & _GEN_3977) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_57_line_3 <= _GEN_2946;
        end else begin
          cache_57_line_3 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_57_line_3 <= _GEN_2169;
      end
    end else begin
      cache_57_line_3 <= _GEN_2169;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_57_line_4 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4882 & _GEN_3979) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_57_line_4 <= _GEN_2946;
        end else begin
          cache_57_line_4 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_57_line_4 <= _GEN_2233;
      end
    end else begin
      cache_57_line_4 <= _GEN_2233;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_57_line_5 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4882 & _GEN_3981) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_57_line_5 <= _GEN_2946;
        end else begin
          cache_57_line_5 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_57_line_5 <= _GEN_2297;
      end
    end else begin
      cache_57_line_5 <= _GEN_2297;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_57_line_6 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4882 & _GEN_3983) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_57_line_6 <= _GEN_2946;
        end else begin
          cache_57_line_6 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_57_line_6 <= _GEN_2361;
      end
    end else begin
      cache_57_line_6 <= _GEN_2361;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_57_line_7 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4882 & _GEN_3985) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_57_line_7 <= _GEN_2946;
        end else begin
          cache_57_line_7 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_57_line_7 <= _GEN_2425;
      end
    end else begin
      cache_57_line_7 <= _GEN_2425;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_58_validBit <= 1'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      cache_58_validBit <= _GEN_1210;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_58_tag <= 5'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      if (6'h3a == cacheLine) begin // @[Cache.scala 50:26]
        cache_58_tag <= tag; // @[Cache.scala 50:26]
      end
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_58_line_0 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4898 & _GEN_3987) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_58_line_0 <= _GEN_2946;
        end else begin
          cache_58_line_0 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_58_line_0 <= _GEN_1978;
      end
    end else begin
      cache_58_line_0 <= _GEN_1978;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_58_line_1 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4898 & _GEN_3973) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_58_line_1 <= _GEN_2946;
        end else begin
          cache_58_line_1 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_58_line_1 <= _GEN_2042;
      end
    end else begin
      cache_58_line_1 <= _GEN_2042;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_58_line_2 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4898 & _GEN_3975) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_58_line_2 <= _GEN_2946;
        end else begin
          cache_58_line_2 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_58_line_2 <= _GEN_2106;
      end
    end else begin
      cache_58_line_2 <= _GEN_2106;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_58_line_3 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4898 & _GEN_3977) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_58_line_3 <= _GEN_2946;
        end else begin
          cache_58_line_3 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_58_line_3 <= _GEN_2170;
      end
    end else begin
      cache_58_line_3 <= _GEN_2170;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_58_line_4 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4898 & _GEN_3979) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_58_line_4 <= _GEN_2946;
        end else begin
          cache_58_line_4 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_58_line_4 <= _GEN_2234;
      end
    end else begin
      cache_58_line_4 <= _GEN_2234;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_58_line_5 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4898 & _GEN_3981) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_58_line_5 <= _GEN_2946;
        end else begin
          cache_58_line_5 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_58_line_5 <= _GEN_2298;
      end
    end else begin
      cache_58_line_5 <= _GEN_2298;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_58_line_6 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4898 & _GEN_3983) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_58_line_6 <= _GEN_2946;
        end else begin
          cache_58_line_6 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_58_line_6 <= _GEN_2362;
      end
    end else begin
      cache_58_line_6 <= _GEN_2362;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_58_line_7 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4898 & _GEN_3985) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_58_line_7 <= _GEN_2946;
        end else begin
          cache_58_line_7 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_58_line_7 <= _GEN_2426;
      end
    end else begin
      cache_58_line_7 <= _GEN_2426;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_59_validBit <= 1'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      cache_59_validBit <= _GEN_1211;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_59_tag <= 5'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      if (6'h3b == cacheLine) begin // @[Cache.scala 50:26]
        cache_59_tag <= tag; // @[Cache.scala 50:26]
      end
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_59_line_0 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4914 & _GEN_3987) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_59_line_0 <= _GEN_2946;
        end else begin
          cache_59_line_0 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_59_line_0 <= _GEN_1979;
      end
    end else begin
      cache_59_line_0 <= _GEN_1979;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_59_line_1 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4914 & _GEN_3973) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_59_line_1 <= _GEN_2946;
        end else begin
          cache_59_line_1 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_59_line_1 <= _GEN_2043;
      end
    end else begin
      cache_59_line_1 <= _GEN_2043;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_59_line_2 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4914 & _GEN_3975) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_59_line_2 <= _GEN_2946;
        end else begin
          cache_59_line_2 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_59_line_2 <= _GEN_2107;
      end
    end else begin
      cache_59_line_2 <= _GEN_2107;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_59_line_3 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4914 & _GEN_3977) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_59_line_3 <= _GEN_2946;
        end else begin
          cache_59_line_3 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_59_line_3 <= _GEN_2171;
      end
    end else begin
      cache_59_line_3 <= _GEN_2171;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_59_line_4 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4914 & _GEN_3979) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_59_line_4 <= _GEN_2946;
        end else begin
          cache_59_line_4 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_59_line_4 <= _GEN_2235;
      end
    end else begin
      cache_59_line_4 <= _GEN_2235;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_59_line_5 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4914 & _GEN_3981) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_59_line_5 <= _GEN_2946;
        end else begin
          cache_59_line_5 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_59_line_5 <= _GEN_2299;
      end
    end else begin
      cache_59_line_5 <= _GEN_2299;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_59_line_6 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4914 & _GEN_3983) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_59_line_6 <= _GEN_2946;
        end else begin
          cache_59_line_6 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_59_line_6 <= _GEN_2363;
      end
    end else begin
      cache_59_line_6 <= _GEN_2363;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_59_line_7 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4914 & _GEN_3985) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_59_line_7 <= _GEN_2946;
        end else begin
          cache_59_line_7 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_59_line_7 <= _GEN_2427;
      end
    end else begin
      cache_59_line_7 <= _GEN_2427;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_60_validBit <= 1'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      cache_60_validBit <= _GEN_1212;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_60_tag <= 5'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      if (6'h3c == cacheLine) begin // @[Cache.scala 50:26]
        cache_60_tag <= tag; // @[Cache.scala 50:26]
      end
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_60_line_0 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4930 & _GEN_3987) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_60_line_0 <= _GEN_2946;
        end else begin
          cache_60_line_0 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_60_line_0 <= _GEN_1980;
      end
    end else begin
      cache_60_line_0 <= _GEN_1980;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_60_line_1 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4930 & _GEN_3973) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_60_line_1 <= _GEN_2946;
        end else begin
          cache_60_line_1 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_60_line_1 <= _GEN_2044;
      end
    end else begin
      cache_60_line_1 <= _GEN_2044;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_60_line_2 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4930 & _GEN_3975) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_60_line_2 <= _GEN_2946;
        end else begin
          cache_60_line_2 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_60_line_2 <= _GEN_2108;
      end
    end else begin
      cache_60_line_2 <= _GEN_2108;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_60_line_3 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4930 & _GEN_3977) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_60_line_3 <= _GEN_2946;
        end else begin
          cache_60_line_3 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_60_line_3 <= _GEN_2172;
      end
    end else begin
      cache_60_line_3 <= _GEN_2172;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_60_line_4 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4930 & _GEN_3979) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_60_line_4 <= _GEN_2946;
        end else begin
          cache_60_line_4 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_60_line_4 <= _GEN_2236;
      end
    end else begin
      cache_60_line_4 <= _GEN_2236;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_60_line_5 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4930 & _GEN_3981) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_60_line_5 <= _GEN_2946;
        end else begin
          cache_60_line_5 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_60_line_5 <= _GEN_2300;
      end
    end else begin
      cache_60_line_5 <= _GEN_2300;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_60_line_6 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4930 & _GEN_3983) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_60_line_6 <= _GEN_2946;
        end else begin
          cache_60_line_6 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_60_line_6 <= _GEN_2364;
      end
    end else begin
      cache_60_line_6 <= _GEN_2364;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_60_line_7 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4930 & _GEN_3985) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_60_line_7 <= _GEN_2946;
        end else begin
          cache_60_line_7 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_60_line_7 <= _GEN_2428;
      end
    end else begin
      cache_60_line_7 <= _GEN_2428;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_61_validBit <= 1'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      cache_61_validBit <= _GEN_1213;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_61_tag <= 5'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      if (6'h3d == cacheLine) begin // @[Cache.scala 50:26]
        cache_61_tag <= tag; // @[Cache.scala 50:26]
      end
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_61_line_0 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4946 & _GEN_3987) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_61_line_0 <= _GEN_2946;
        end else begin
          cache_61_line_0 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_61_line_0 <= _GEN_1981;
      end
    end else begin
      cache_61_line_0 <= _GEN_1981;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_61_line_1 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4946 & _GEN_3973) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_61_line_1 <= _GEN_2946;
        end else begin
          cache_61_line_1 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_61_line_1 <= _GEN_2045;
      end
    end else begin
      cache_61_line_1 <= _GEN_2045;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_61_line_2 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4946 & _GEN_3975) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_61_line_2 <= _GEN_2946;
        end else begin
          cache_61_line_2 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_61_line_2 <= _GEN_2109;
      end
    end else begin
      cache_61_line_2 <= _GEN_2109;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_61_line_3 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4946 & _GEN_3977) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_61_line_3 <= _GEN_2946;
        end else begin
          cache_61_line_3 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_61_line_3 <= _GEN_2173;
      end
    end else begin
      cache_61_line_3 <= _GEN_2173;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_61_line_4 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4946 & _GEN_3979) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_61_line_4 <= _GEN_2946;
        end else begin
          cache_61_line_4 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_61_line_4 <= _GEN_2237;
      end
    end else begin
      cache_61_line_4 <= _GEN_2237;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_61_line_5 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4946 & _GEN_3981) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_61_line_5 <= _GEN_2946;
        end else begin
          cache_61_line_5 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_61_line_5 <= _GEN_2301;
      end
    end else begin
      cache_61_line_5 <= _GEN_2301;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_61_line_6 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4946 & _GEN_3983) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_61_line_6 <= _GEN_2946;
        end else begin
          cache_61_line_6 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_61_line_6 <= _GEN_2365;
      end
    end else begin
      cache_61_line_6 <= _GEN_2365;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_61_line_7 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4946 & _GEN_3985) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_61_line_7 <= _GEN_2946;
        end else begin
          cache_61_line_7 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_61_line_7 <= _GEN_2429;
      end
    end else begin
      cache_61_line_7 <= _GEN_2429;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_62_validBit <= 1'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      cache_62_validBit <= _GEN_1214;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_62_tag <= 5'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      if (6'h3e == cacheLine) begin // @[Cache.scala 50:26]
        cache_62_tag <= tag; // @[Cache.scala 50:26]
      end
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_62_line_0 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4962 & _GEN_3987) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_62_line_0 <= _GEN_2946;
        end else begin
          cache_62_line_0 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_62_line_0 <= _GEN_1982;
      end
    end else begin
      cache_62_line_0 <= _GEN_1982;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_62_line_1 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4962 & _GEN_3973) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_62_line_1 <= _GEN_2946;
        end else begin
          cache_62_line_1 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_62_line_1 <= _GEN_2046;
      end
    end else begin
      cache_62_line_1 <= _GEN_2046;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_62_line_2 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4962 & _GEN_3975) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_62_line_2 <= _GEN_2946;
        end else begin
          cache_62_line_2 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_62_line_2 <= _GEN_2110;
      end
    end else begin
      cache_62_line_2 <= _GEN_2110;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_62_line_3 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4962 & _GEN_3977) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_62_line_3 <= _GEN_2946;
        end else begin
          cache_62_line_3 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_62_line_3 <= _GEN_2174;
      end
    end else begin
      cache_62_line_3 <= _GEN_2174;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_62_line_4 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4962 & _GEN_3979) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_62_line_4 <= _GEN_2946;
        end else begin
          cache_62_line_4 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_62_line_4 <= _GEN_2238;
      end
    end else begin
      cache_62_line_4 <= _GEN_2238;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_62_line_5 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4962 & _GEN_3981) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_62_line_5 <= _GEN_2946;
        end else begin
          cache_62_line_5 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_62_line_5 <= _GEN_2302;
      end
    end else begin
      cache_62_line_5 <= _GEN_2302;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_62_line_6 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4962 & _GEN_3983) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_62_line_6 <= _GEN_2946;
        end else begin
          cache_62_line_6 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_62_line_6 <= _GEN_2366;
      end
    end else begin
      cache_62_line_6 <= _GEN_2366;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_62_line_7 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4962 & _GEN_3985) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_62_line_7 <= _GEN_2946;
        end else begin
          cache_62_line_7 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_62_line_7 <= _GEN_2430;
      end
    end else begin
      cache_62_line_7 <= _GEN_2430;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_63_validBit <= 1'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      cache_63_validBit <= _GEN_1215;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_63_tag <= 5'h0; // @[Cache.scala 32:22]
    end else if (io_blockWriteEn) begin // @[Cache.scala 48:25]
      if (6'h3f == cacheLine) begin // @[Cache.scala 50:26]
        cache_63_tag <= tag; // @[Cache.scala 50:26]
      end
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_63_line_0 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4978 & _GEN_3987) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_63_line_0 <= _GEN_2946;
        end else begin
          cache_63_line_0 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_63_line_0 <= _GEN_1983;
      end
    end else begin
      cache_63_line_0 <= _GEN_1983;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_63_line_1 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4978 & _GEN_3973) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_63_line_1 <= _GEN_2946;
        end else begin
          cache_63_line_1 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_63_line_1 <= _GEN_2047;
      end
    end else begin
      cache_63_line_1 <= _GEN_2047;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_63_line_2 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4978 & _GEN_3975) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_63_line_2 <= _GEN_2946;
        end else begin
          cache_63_line_2 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_63_line_2 <= _GEN_2111;
      end
    end else begin
      cache_63_line_2 <= _GEN_2111;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_63_line_3 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4978 & _GEN_3977) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_63_line_3 <= _GEN_2946;
        end else begin
          cache_63_line_3 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_63_line_3 <= _GEN_2175;
      end
    end else begin
      cache_63_line_3 <= _GEN_2175;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_63_line_4 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4978 & _GEN_3979) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_63_line_4 <= _GEN_2946;
        end else begin
          cache_63_line_4 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_63_line_4 <= _GEN_2239;
      end
    end else begin
      cache_63_line_4 <= _GEN_2239;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_63_line_5 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4978 & _GEN_3981) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_63_line_5 <= _GEN_2946;
        end else begin
          cache_63_line_5 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_63_line_5 <= _GEN_2303;
      end
    end else begin
      cache_63_line_5 <= _GEN_2303;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_63_line_6 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4978 & _GEN_3983) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_63_line_6 <= _GEN_2946;
        end else begin
          cache_63_line_6 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_63_line_6 <= _GEN_2367;
      end
    end else begin
      cache_63_line_6 <= _GEN_2367;
    end
    if (reset) begin // @[Cache.scala 32:22]
      cache_63_line_7 <= 32'h0; // @[Cache.scala 32:22]
    end else if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
      if (_GEN_4978 & _GEN_3985) begin // @[Cache.scala 71:43]
        if (io_cpuWriteEn & hit) begin // @[Cache.scala 59:29]
          cache_63_line_7 <= _GEN_2946;
        end else begin
          cache_63_line_7 <= 32'h0; // @[Cache.scala 57:30]
        end
      end else begin
        cache_63_line_7 <= _GEN_2431;
      end
    end else begin
      cache_63_line_7 <= _GEN_2431;
    end
    if (reset) begin // @[Cache.scala 33:27]
      dataBuffer <= 256'h0; // @[Cache.scala 33:27]
    end else begin
      dataBuffer <= _dataBuffer_T; // @[Cache.scala 45:14]
    end
    if (reset) begin // @[Cache.scala 34:28]
      addrsBuffer <= 16'h0; // @[Cache.scala 34:28]
    end else begin
      addrsBuffer <= {{5'd0}, _addrsBuffer_T}; // @[Cache.scala 44:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cache_0_validBit = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  cache_0_tag = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  cache_0_line_0 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  cache_0_line_1 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  cache_0_line_2 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  cache_0_line_3 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  cache_0_line_4 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  cache_0_line_5 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  cache_0_line_6 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  cache_0_line_7 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  cache_1_validBit = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  cache_1_tag = _RAND_11[4:0];
  _RAND_12 = {1{`RANDOM}};
  cache_1_line_0 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  cache_1_line_1 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  cache_1_line_2 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  cache_1_line_3 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  cache_1_line_4 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  cache_1_line_5 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  cache_1_line_6 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  cache_1_line_7 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  cache_2_validBit = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  cache_2_tag = _RAND_21[4:0];
  _RAND_22 = {1{`RANDOM}};
  cache_2_line_0 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  cache_2_line_1 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  cache_2_line_2 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  cache_2_line_3 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  cache_2_line_4 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  cache_2_line_5 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  cache_2_line_6 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  cache_2_line_7 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  cache_3_validBit = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  cache_3_tag = _RAND_31[4:0];
  _RAND_32 = {1{`RANDOM}};
  cache_3_line_0 = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  cache_3_line_1 = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  cache_3_line_2 = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  cache_3_line_3 = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  cache_3_line_4 = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  cache_3_line_5 = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  cache_3_line_6 = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  cache_3_line_7 = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  cache_4_validBit = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  cache_4_tag = _RAND_41[4:0];
  _RAND_42 = {1{`RANDOM}};
  cache_4_line_0 = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  cache_4_line_1 = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  cache_4_line_2 = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  cache_4_line_3 = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  cache_4_line_4 = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  cache_4_line_5 = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  cache_4_line_6 = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  cache_4_line_7 = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  cache_5_validBit = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  cache_5_tag = _RAND_51[4:0];
  _RAND_52 = {1{`RANDOM}};
  cache_5_line_0 = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  cache_5_line_1 = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  cache_5_line_2 = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  cache_5_line_3 = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  cache_5_line_4 = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  cache_5_line_5 = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  cache_5_line_6 = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  cache_5_line_7 = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  cache_6_validBit = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  cache_6_tag = _RAND_61[4:0];
  _RAND_62 = {1{`RANDOM}};
  cache_6_line_0 = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  cache_6_line_1 = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  cache_6_line_2 = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  cache_6_line_3 = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  cache_6_line_4 = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  cache_6_line_5 = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  cache_6_line_6 = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  cache_6_line_7 = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  cache_7_validBit = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  cache_7_tag = _RAND_71[4:0];
  _RAND_72 = {1{`RANDOM}};
  cache_7_line_0 = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  cache_7_line_1 = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  cache_7_line_2 = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  cache_7_line_3 = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  cache_7_line_4 = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  cache_7_line_5 = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  cache_7_line_6 = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  cache_7_line_7 = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  cache_8_validBit = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  cache_8_tag = _RAND_81[4:0];
  _RAND_82 = {1{`RANDOM}};
  cache_8_line_0 = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  cache_8_line_1 = _RAND_83[31:0];
  _RAND_84 = {1{`RANDOM}};
  cache_8_line_2 = _RAND_84[31:0];
  _RAND_85 = {1{`RANDOM}};
  cache_8_line_3 = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  cache_8_line_4 = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  cache_8_line_5 = _RAND_87[31:0];
  _RAND_88 = {1{`RANDOM}};
  cache_8_line_6 = _RAND_88[31:0];
  _RAND_89 = {1{`RANDOM}};
  cache_8_line_7 = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  cache_9_validBit = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  cache_9_tag = _RAND_91[4:0];
  _RAND_92 = {1{`RANDOM}};
  cache_9_line_0 = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  cache_9_line_1 = _RAND_93[31:0];
  _RAND_94 = {1{`RANDOM}};
  cache_9_line_2 = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  cache_9_line_3 = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  cache_9_line_4 = _RAND_96[31:0];
  _RAND_97 = {1{`RANDOM}};
  cache_9_line_5 = _RAND_97[31:0];
  _RAND_98 = {1{`RANDOM}};
  cache_9_line_6 = _RAND_98[31:0];
  _RAND_99 = {1{`RANDOM}};
  cache_9_line_7 = _RAND_99[31:0];
  _RAND_100 = {1{`RANDOM}};
  cache_10_validBit = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  cache_10_tag = _RAND_101[4:0];
  _RAND_102 = {1{`RANDOM}};
  cache_10_line_0 = _RAND_102[31:0];
  _RAND_103 = {1{`RANDOM}};
  cache_10_line_1 = _RAND_103[31:0];
  _RAND_104 = {1{`RANDOM}};
  cache_10_line_2 = _RAND_104[31:0];
  _RAND_105 = {1{`RANDOM}};
  cache_10_line_3 = _RAND_105[31:0];
  _RAND_106 = {1{`RANDOM}};
  cache_10_line_4 = _RAND_106[31:0];
  _RAND_107 = {1{`RANDOM}};
  cache_10_line_5 = _RAND_107[31:0];
  _RAND_108 = {1{`RANDOM}};
  cache_10_line_6 = _RAND_108[31:0];
  _RAND_109 = {1{`RANDOM}};
  cache_10_line_7 = _RAND_109[31:0];
  _RAND_110 = {1{`RANDOM}};
  cache_11_validBit = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  cache_11_tag = _RAND_111[4:0];
  _RAND_112 = {1{`RANDOM}};
  cache_11_line_0 = _RAND_112[31:0];
  _RAND_113 = {1{`RANDOM}};
  cache_11_line_1 = _RAND_113[31:0];
  _RAND_114 = {1{`RANDOM}};
  cache_11_line_2 = _RAND_114[31:0];
  _RAND_115 = {1{`RANDOM}};
  cache_11_line_3 = _RAND_115[31:0];
  _RAND_116 = {1{`RANDOM}};
  cache_11_line_4 = _RAND_116[31:0];
  _RAND_117 = {1{`RANDOM}};
  cache_11_line_5 = _RAND_117[31:0];
  _RAND_118 = {1{`RANDOM}};
  cache_11_line_6 = _RAND_118[31:0];
  _RAND_119 = {1{`RANDOM}};
  cache_11_line_7 = _RAND_119[31:0];
  _RAND_120 = {1{`RANDOM}};
  cache_12_validBit = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  cache_12_tag = _RAND_121[4:0];
  _RAND_122 = {1{`RANDOM}};
  cache_12_line_0 = _RAND_122[31:0];
  _RAND_123 = {1{`RANDOM}};
  cache_12_line_1 = _RAND_123[31:0];
  _RAND_124 = {1{`RANDOM}};
  cache_12_line_2 = _RAND_124[31:0];
  _RAND_125 = {1{`RANDOM}};
  cache_12_line_3 = _RAND_125[31:0];
  _RAND_126 = {1{`RANDOM}};
  cache_12_line_4 = _RAND_126[31:0];
  _RAND_127 = {1{`RANDOM}};
  cache_12_line_5 = _RAND_127[31:0];
  _RAND_128 = {1{`RANDOM}};
  cache_12_line_6 = _RAND_128[31:0];
  _RAND_129 = {1{`RANDOM}};
  cache_12_line_7 = _RAND_129[31:0];
  _RAND_130 = {1{`RANDOM}};
  cache_13_validBit = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  cache_13_tag = _RAND_131[4:0];
  _RAND_132 = {1{`RANDOM}};
  cache_13_line_0 = _RAND_132[31:0];
  _RAND_133 = {1{`RANDOM}};
  cache_13_line_1 = _RAND_133[31:0];
  _RAND_134 = {1{`RANDOM}};
  cache_13_line_2 = _RAND_134[31:0];
  _RAND_135 = {1{`RANDOM}};
  cache_13_line_3 = _RAND_135[31:0];
  _RAND_136 = {1{`RANDOM}};
  cache_13_line_4 = _RAND_136[31:0];
  _RAND_137 = {1{`RANDOM}};
  cache_13_line_5 = _RAND_137[31:0];
  _RAND_138 = {1{`RANDOM}};
  cache_13_line_6 = _RAND_138[31:0];
  _RAND_139 = {1{`RANDOM}};
  cache_13_line_7 = _RAND_139[31:0];
  _RAND_140 = {1{`RANDOM}};
  cache_14_validBit = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  cache_14_tag = _RAND_141[4:0];
  _RAND_142 = {1{`RANDOM}};
  cache_14_line_0 = _RAND_142[31:0];
  _RAND_143 = {1{`RANDOM}};
  cache_14_line_1 = _RAND_143[31:0];
  _RAND_144 = {1{`RANDOM}};
  cache_14_line_2 = _RAND_144[31:0];
  _RAND_145 = {1{`RANDOM}};
  cache_14_line_3 = _RAND_145[31:0];
  _RAND_146 = {1{`RANDOM}};
  cache_14_line_4 = _RAND_146[31:0];
  _RAND_147 = {1{`RANDOM}};
  cache_14_line_5 = _RAND_147[31:0];
  _RAND_148 = {1{`RANDOM}};
  cache_14_line_6 = _RAND_148[31:0];
  _RAND_149 = {1{`RANDOM}};
  cache_14_line_7 = _RAND_149[31:0];
  _RAND_150 = {1{`RANDOM}};
  cache_15_validBit = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  cache_15_tag = _RAND_151[4:0];
  _RAND_152 = {1{`RANDOM}};
  cache_15_line_0 = _RAND_152[31:0];
  _RAND_153 = {1{`RANDOM}};
  cache_15_line_1 = _RAND_153[31:0];
  _RAND_154 = {1{`RANDOM}};
  cache_15_line_2 = _RAND_154[31:0];
  _RAND_155 = {1{`RANDOM}};
  cache_15_line_3 = _RAND_155[31:0];
  _RAND_156 = {1{`RANDOM}};
  cache_15_line_4 = _RAND_156[31:0];
  _RAND_157 = {1{`RANDOM}};
  cache_15_line_5 = _RAND_157[31:0];
  _RAND_158 = {1{`RANDOM}};
  cache_15_line_6 = _RAND_158[31:0];
  _RAND_159 = {1{`RANDOM}};
  cache_15_line_7 = _RAND_159[31:0];
  _RAND_160 = {1{`RANDOM}};
  cache_16_validBit = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  cache_16_tag = _RAND_161[4:0];
  _RAND_162 = {1{`RANDOM}};
  cache_16_line_0 = _RAND_162[31:0];
  _RAND_163 = {1{`RANDOM}};
  cache_16_line_1 = _RAND_163[31:0];
  _RAND_164 = {1{`RANDOM}};
  cache_16_line_2 = _RAND_164[31:0];
  _RAND_165 = {1{`RANDOM}};
  cache_16_line_3 = _RAND_165[31:0];
  _RAND_166 = {1{`RANDOM}};
  cache_16_line_4 = _RAND_166[31:0];
  _RAND_167 = {1{`RANDOM}};
  cache_16_line_5 = _RAND_167[31:0];
  _RAND_168 = {1{`RANDOM}};
  cache_16_line_6 = _RAND_168[31:0];
  _RAND_169 = {1{`RANDOM}};
  cache_16_line_7 = _RAND_169[31:0];
  _RAND_170 = {1{`RANDOM}};
  cache_17_validBit = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  cache_17_tag = _RAND_171[4:0];
  _RAND_172 = {1{`RANDOM}};
  cache_17_line_0 = _RAND_172[31:0];
  _RAND_173 = {1{`RANDOM}};
  cache_17_line_1 = _RAND_173[31:0];
  _RAND_174 = {1{`RANDOM}};
  cache_17_line_2 = _RAND_174[31:0];
  _RAND_175 = {1{`RANDOM}};
  cache_17_line_3 = _RAND_175[31:0];
  _RAND_176 = {1{`RANDOM}};
  cache_17_line_4 = _RAND_176[31:0];
  _RAND_177 = {1{`RANDOM}};
  cache_17_line_5 = _RAND_177[31:0];
  _RAND_178 = {1{`RANDOM}};
  cache_17_line_6 = _RAND_178[31:0];
  _RAND_179 = {1{`RANDOM}};
  cache_17_line_7 = _RAND_179[31:0];
  _RAND_180 = {1{`RANDOM}};
  cache_18_validBit = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  cache_18_tag = _RAND_181[4:0];
  _RAND_182 = {1{`RANDOM}};
  cache_18_line_0 = _RAND_182[31:0];
  _RAND_183 = {1{`RANDOM}};
  cache_18_line_1 = _RAND_183[31:0];
  _RAND_184 = {1{`RANDOM}};
  cache_18_line_2 = _RAND_184[31:0];
  _RAND_185 = {1{`RANDOM}};
  cache_18_line_3 = _RAND_185[31:0];
  _RAND_186 = {1{`RANDOM}};
  cache_18_line_4 = _RAND_186[31:0];
  _RAND_187 = {1{`RANDOM}};
  cache_18_line_5 = _RAND_187[31:0];
  _RAND_188 = {1{`RANDOM}};
  cache_18_line_6 = _RAND_188[31:0];
  _RAND_189 = {1{`RANDOM}};
  cache_18_line_7 = _RAND_189[31:0];
  _RAND_190 = {1{`RANDOM}};
  cache_19_validBit = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  cache_19_tag = _RAND_191[4:0];
  _RAND_192 = {1{`RANDOM}};
  cache_19_line_0 = _RAND_192[31:0];
  _RAND_193 = {1{`RANDOM}};
  cache_19_line_1 = _RAND_193[31:0];
  _RAND_194 = {1{`RANDOM}};
  cache_19_line_2 = _RAND_194[31:0];
  _RAND_195 = {1{`RANDOM}};
  cache_19_line_3 = _RAND_195[31:0];
  _RAND_196 = {1{`RANDOM}};
  cache_19_line_4 = _RAND_196[31:0];
  _RAND_197 = {1{`RANDOM}};
  cache_19_line_5 = _RAND_197[31:0];
  _RAND_198 = {1{`RANDOM}};
  cache_19_line_6 = _RAND_198[31:0];
  _RAND_199 = {1{`RANDOM}};
  cache_19_line_7 = _RAND_199[31:0];
  _RAND_200 = {1{`RANDOM}};
  cache_20_validBit = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  cache_20_tag = _RAND_201[4:0];
  _RAND_202 = {1{`RANDOM}};
  cache_20_line_0 = _RAND_202[31:0];
  _RAND_203 = {1{`RANDOM}};
  cache_20_line_1 = _RAND_203[31:0];
  _RAND_204 = {1{`RANDOM}};
  cache_20_line_2 = _RAND_204[31:0];
  _RAND_205 = {1{`RANDOM}};
  cache_20_line_3 = _RAND_205[31:0];
  _RAND_206 = {1{`RANDOM}};
  cache_20_line_4 = _RAND_206[31:0];
  _RAND_207 = {1{`RANDOM}};
  cache_20_line_5 = _RAND_207[31:0];
  _RAND_208 = {1{`RANDOM}};
  cache_20_line_6 = _RAND_208[31:0];
  _RAND_209 = {1{`RANDOM}};
  cache_20_line_7 = _RAND_209[31:0];
  _RAND_210 = {1{`RANDOM}};
  cache_21_validBit = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  cache_21_tag = _RAND_211[4:0];
  _RAND_212 = {1{`RANDOM}};
  cache_21_line_0 = _RAND_212[31:0];
  _RAND_213 = {1{`RANDOM}};
  cache_21_line_1 = _RAND_213[31:0];
  _RAND_214 = {1{`RANDOM}};
  cache_21_line_2 = _RAND_214[31:0];
  _RAND_215 = {1{`RANDOM}};
  cache_21_line_3 = _RAND_215[31:0];
  _RAND_216 = {1{`RANDOM}};
  cache_21_line_4 = _RAND_216[31:0];
  _RAND_217 = {1{`RANDOM}};
  cache_21_line_5 = _RAND_217[31:0];
  _RAND_218 = {1{`RANDOM}};
  cache_21_line_6 = _RAND_218[31:0];
  _RAND_219 = {1{`RANDOM}};
  cache_21_line_7 = _RAND_219[31:0];
  _RAND_220 = {1{`RANDOM}};
  cache_22_validBit = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  cache_22_tag = _RAND_221[4:0];
  _RAND_222 = {1{`RANDOM}};
  cache_22_line_0 = _RAND_222[31:0];
  _RAND_223 = {1{`RANDOM}};
  cache_22_line_1 = _RAND_223[31:0];
  _RAND_224 = {1{`RANDOM}};
  cache_22_line_2 = _RAND_224[31:0];
  _RAND_225 = {1{`RANDOM}};
  cache_22_line_3 = _RAND_225[31:0];
  _RAND_226 = {1{`RANDOM}};
  cache_22_line_4 = _RAND_226[31:0];
  _RAND_227 = {1{`RANDOM}};
  cache_22_line_5 = _RAND_227[31:0];
  _RAND_228 = {1{`RANDOM}};
  cache_22_line_6 = _RAND_228[31:0];
  _RAND_229 = {1{`RANDOM}};
  cache_22_line_7 = _RAND_229[31:0];
  _RAND_230 = {1{`RANDOM}};
  cache_23_validBit = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  cache_23_tag = _RAND_231[4:0];
  _RAND_232 = {1{`RANDOM}};
  cache_23_line_0 = _RAND_232[31:0];
  _RAND_233 = {1{`RANDOM}};
  cache_23_line_1 = _RAND_233[31:0];
  _RAND_234 = {1{`RANDOM}};
  cache_23_line_2 = _RAND_234[31:0];
  _RAND_235 = {1{`RANDOM}};
  cache_23_line_3 = _RAND_235[31:0];
  _RAND_236 = {1{`RANDOM}};
  cache_23_line_4 = _RAND_236[31:0];
  _RAND_237 = {1{`RANDOM}};
  cache_23_line_5 = _RAND_237[31:0];
  _RAND_238 = {1{`RANDOM}};
  cache_23_line_6 = _RAND_238[31:0];
  _RAND_239 = {1{`RANDOM}};
  cache_23_line_7 = _RAND_239[31:0];
  _RAND_240 = {1{`RANDOM}};
  cache_24_validBit = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  cache_24_tag = _RAND_241[4:0];
  _RAND_242 = {1{`RANDOM}};
  cache_24_line_0 = _RAND_242[31:0];
  _RAND_243 = {1{`RANDOM}};
  cache_24_line_1 = _RAND_243[31:0];
  _RAND_244 = {1{`RANDOM}};
  cache_24_line_2 = _RAND_244[31:0];
  _RAND_245 = {1{`RANDOM}};
  cache_24_line_3 = _RAND_245[31:0];
  _RAND_246 = {1{`RANDOM}};
  cache_24_line_4 = _RAND_246[31:0];
  _RAND_247 = {1{`RANDOM}};
  cache_24_line_5 = _RAND_247[31:0];
  _RAND_248 = {1{`RANDOM}};
  cache_24_line_6 = _RAND_248[31:0];
  _RAND_249 = {1{`RANDOM}};
  cache_24_line_7 = _RAND_249[31:0];
  _RAND_250 = {1{`RANDOM}};
  cache_25_validBit = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  cache_25_tag = _RAND_251[4:0];
  _RAND_252 = {1{`RANDOM}};
  cache_25_line_0 = _RAND_252[31:0];
  _RAND_253 = {1{`RANDOM}};
  cache_25_line_1 = _RAND_253[31:0];
  _RAND_254 = {1{`RANDOM}};
  cache_25_line_2 = _RAND_254[31:0];
  _RAND_255 = {1{`RANDOM}};
  cache_25_line_3 = _RAND_255[31:0];
  _RAND_256 = {1{`RANDOM}};
  cache_25_line_4 = _RAND_256[31:0];
  _RAND_257 = {1{`RANDOM}};
  cache_25_line_5 = _RAND_257[31:0];
  _RAND_258 = {1{`RANDOM}};
  cache_25_line_6 = _RAND_258[31:0];
  _RAND_259 = {1{`RANDOM}};
  cache_25_line_7 = _RAND_259[31:0];
  _RAND_260 = {1{`RANDOM}};
  cache_26_validBit = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  cache_26_tag = _RAND_261[4:0];
  _RAND_262 = {1{`RANDOM}};
  cache_26_line_0 = _RAND_262[31:0];
  _RAND_263 = {1{`RANDOM}};
  cache_26_line_1 = _RAND_263[31:0];
  _RAND_264 = {1{`RANDOM}};
  cache_26_line_2 = _RAND_264[31:0];
  _RAND_265 = {1{`RANDOM}};
  cache_26_line_3 = _RAND_265[31:0];
  _RAND_266 = {1{`RANDOM}};
  cache_26_line_4 = _RAND_266[31:0];
  _RAND_267 = {1{`RANDOM}};
  cache_26_line_5 = _RAND_267[31:0];
  _RAND_268 = {1{`RANDOM}};
  cache_26_line_6 = _RAND_268[31:0];
  _RAND_269 = {1{`RANDOM}};
  cache_26_line_7 = _RAND_269[31:0];
  _RAND_270 = {1{`RANDOM}};
  cache_27_validBit = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  cache_27_tag = _RAND_271[4:0];
  _RAND_272 = {1{`RANDOM}};
  cache_27_line_0 = _RAND_272[31:0];
  _RAND_273 = {1{`RANDOM}};
  cache_27_line_1 = _RAND_273[31:0];
  _RAND_274 = {1{`RANDOM}};
  cache_27_line_2 = _RAND_274[31:0];
  _RAND_275 = {1{`RANDOM}};
  cache_27_line_3 = _RAND_275[31:0];
  _RAND_276 = {1{`RANDOM}};
  cache_27_line_4 = _RAND_276[31:0];
  _RAND_277 = {1{`RANDOM}};
  cache_27_line_5 = _RAND_277[31:0];
  _RAND_278 = {1{`RANDOM}};
  cache_27_line_6 = _RAND_278[31:0];
  _RAND_279 = {1{`RANDOM}};
  cache_27_line_7 = _RAND_279[31:0];
  _RAND_280 = {1{`RANDOM}};
  cache_28_validBit = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  cache_28_tag = _RAND_281[4:0];
  _RAND_282 = {1{`RANDOM}};
  cache_28_line_0 = _RAND_282[31:0];
  _RAND_283 = {1{`RANDOM}};
  cache_28_line_1 = _RAND_283[31:0];
  _RAND_284 = {1{`RANDOM}};
  cache_28_line_2 = _RAND_284[31:0];
  _RAND_285 = {1{`RANDOM}};
  cache_28_line_3 = _RAND_285[31:0];
  _RAND_286 = {1{`RANDOM}};
  cache_28_line_4 = _RAND_286[31:0];
  _RAND_287 = {1{`RANDOM}};
  cache_28_line_5 = _RAND_287[31:0];
  _RAND_288 = {1{`RANDOM}};
  cache_28_line_6 = _RAND_288[31:0];
  _RAND_289 = {1{`RANDOM}};
  cache_28_line_7 = _RAND_289[31:0];
  _RAND_290 = {1{`RANDOM}};
  cache_29_validBit = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  cache_29_tag = _RAND_291[4:0];
  _RAND_292 = {1{`RANDOM}};
  cache_29_line_0 = _RAND_292[31:0];
  _RAND_293 = {1{`RANDOM}};
  cache_29_line_1 = _RAND_293[31:0];
  _RAND_294 = {1{`RANDOM}};
  cache_29_line_2 = _RAND_294[31:0];
  _RAND_295 = {1{`RANDOM}};
  cache_29_line_3 = _RAND_295[31:0];
  _RAND_296 = {1{`RANDOM}};
  cache_29_line_4 = _RAND_296[31:0];
  _RAND_297 = {1{`RANDOM}};
  cache_29_line_5 = _RAND_297[31:0];
  _RAND_298 = {1{`RANDOM}};
  cache_29_line_6 = _RAND_298[31:0];
  _RAND_299 = {1{`RANDOM}};
  cache_29_line_7 = _RAND_299[31:0];
  _RAND_300 = {1{`RANDOM}};
  cache_30_validBit = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  cache_30_tag = _RAND_301[4:0];
  _RAND_302 = {1{`RANDOM}};
  cache_30_line_0 = _RAND_302[31:0];
  _RAND_303 = {1{`RANDOM}};
  cache_30_line_1 = _RAND_303[31:0];
  _RAND_304 = {1{`RANDOM}};
  cache_30_line_2 = _RAND_304[31:0];
  _RAND_305 = {1{`RANDOM}};
  cache_30_line_3 = _RAND_305[31:0];
  _RAND_306 = {1{`RANDOM}};
  cache_30_line_4 = _RAND_306[31:0];
  _RAND_307 = {1{`RANDOM}};
  cache_30_line_5 = _RAND_307[31:0];
  _RAND_308 = {1{`RANDOM}};
  cache_30_line_6 = _RAND_308[31:0];
  _RAND_309 = {1{`RANDOM}};
  cache_30_line_7 = _RAND_309[31:0];
  _RAND_310 = {1{`RANDOM}};
  cache_31_validBit = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  cache_31_tag = _RAND_311[4:0];
  _RAND_312 = {1{`RANDOM}};
  cache_31_line_0 = _RAND_312[31:0];
  _RAND_313 = {1{`RANDOM}};
  cache_31_line_1 = _RAND_313[31:0];
  _RAND_314 = {1{`RANDOM}};
  cache_31_line_2 = _RAND_314[31:0];
  _RAND_315 = {1{`RANDOM}};
  cache_31_line_3 = _RAND_315[31:0];
  _RAND_316 = {1{`RANDOM}};
  cache_31_line_4 = _RAND_316[31:0];
  _RAND_317 = {1{`RANDOM}};
  cache_31_line_5 = _RAND_317[31:0];
  _RAND_318 = {1{`RANDOM}};
  cache_31_line_6 = _RAND_318[31:0];
  _RAND_319 = {1{`RANDOM}};
  cache_31_line_7 = _RAND_319[31:0];
  _RAND_320 = {1{`RANDOM}};
  cache_32_validBit = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  cache_32_tag = _RAND_321[4:0];
  _RAND_322 = {1{`RANDOM}};
  cache_32_line_0 = _RAND_322[31:0];
  _RAND_323 = {1{`RANDOM}};
  cache_32_line_1 = _RAND_323[31:0];
  _RAND_324 = {1{`RANDOM}};
  cache_32_line_2 = _RAND_324[31:0];
  _RAND_325 = {1{`RANDOM}};
  cache_32_line_3 = _RAND_325[31:0];
  _RAND_326 = {1{`RANDOM}};
  cache_32_line_4 = _RAND_326[31:0];
  _RAND_327 = {1{`RANDOM}};
  cache_32_line_5 = _RAND_327[31:0];
  _RAND_328 = {1{`RANDOM}};
  cache_32_line_6 = _RAND_328[31:0];
  _RAND_329 = {1{`RANDOM}};
  cache_32_line_7 = _RAND_329[31:0];
  _RAND_330 = {1{`RANDOM}};
  cache_33_validBit = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  cache_33_tag = _RAND_331[4:0];
  _RAND_332 = {1{`RANDOM}};
  cache_33_line_0 = _RAND_332[31:0];
  _RAND_333 = {1{`RANDOM}};
  cache_33_line_1 = _RAND_333[31:0];
  _RAND_334 = {1{`RANDOM}};
  cache_33_line_2 = _RAND_334[31:0];
  _RAND_335 = {1{`RANDOM}};
  cache_33_line_3 = _RAND_335[31:0];
  _RAND_336 = {1{`RANDOM}};
  cache_33_line_4 = _RAND_336[31:0];
  _RAND_337 = {1{`RANDOM}};
  cache_33_line_5 = _RAND_337[31:0];
  _RAND_338 = {1{`RANDOM}};
  cache_33_line_6 = _RAND_338[31:0];
  _RAND_339 = {1{`RANDOM}};
  cache_33_line_7 = _RAND_339[31:0];
  _RAND_340 = {1{`RANDOM}};
  cache_34_validBit = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  cache_34_tag = _RAND_341[4:0];
  _RAND_342 = {1{`RANDOM}};
  cache_34_line_0 = _RAND_342[31:0];
  _RAND_343 = {1{`RANDOM}};
  cache_34_line_1 = _RAND_343[31:0];
  _RAND_344 = {1{`RANDOM}};
  cache_34_line_2 = _RAND_344[31:0];
  _RAND_345 = {1{`RANDOM}};
  cache_34_line_3 = _RAND_345[31:0];
  _RAND_346 = {1{`RANDOM}};
  cache_34_line_4 = _RAND_346[31:0];
  _RAND_347 = {1{`RANDOM}};
  cache_34_line_5 = _RAND_347[31:0];
  _RAND_348 = {1{`RANDOM}};
  cache_34_line_6 = _RAND_348[31:0];
  _RAND_349 = {1{`RANDOM}};
  cache_34_line_7 = _RAND_349[31:0];
  _RAND_350 = {1{`RANDOM}};
  cache_35_validBit = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  cache_35_tag = _RAND_351[4:0];
  _RAND_352 = {1{`RANDOM}};
  cache_35_line_0 = _RAND_352[31:0];
  _RAND_353 = {1{`RANDOM}};
  cache_35_line_1 = _RAND_353[31:0];
  _RAND_354 = {1{`RANDOM}};
  cache_35_line_2 = _RAND_354[31:0];
  _RAND_355 = {1{`RANDOM}};
  cache_35_line_3 = _RAND_355[31:0];
  _RAND_356 = {1{`RANDOM}};
  cache_35_line_4 = _RAND_356[31:0];
  _RAND_357 = {1{`RANDOM}};
  cache_35_line_5 = _RAND_357[31:0];
  _RAND_358 = {1{`RANDOM}};
  cache_35_line_6 = _RAND_358[31:0];
  _RAND_359 = {1{`RANDOM}};
  cache_35_line_7 = _RAND_359[31:0];
  _RAND_360 = {1{`RANDOM}};
  cache_36_validBit = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  cache_36_tag = _RAND_361[4:0];
  _RAND_362 = {1{`RANDOM}};
  cache_36_line_0 = _RAND_362[31:0];
  _RAND_363 = {1{`RANDOM}};
  cache_36_line_1 = _RAND_363[31:0];
  _RAND_364 = {1{`RANDOM}};
  cache_36_line_2 = _RAND_364[31:0];
  _RAND_365 = {1{`RANDOM}};
  cache_36_line_3 = _RAND_365[31:0];
  _RAND_366 = {1{`RANDOM}};
  cache_36_line_4 = _RAND_366[31:0];
  _RAND_367 = {1{`RANDOM}};
  cache_36_line_5 = _RAND_367[31:0];
  _RAND_368 = {1{`RANDOM}};
  cache_36_line_6 = _RAND_368[31:0];
  _RAND_369 = {1{`RANDOM}};
  cache_36_line_7 = _RAND_369[31:0];
  _RAND_370 = {1{`RANDOM}};
  cache_37_validBit = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  cache_37_tag = _RAND_371[4:0];
  _RAND_372 = {1{`RANDOM}};
  cache_37_line_0 = _RAND_372[31:0];
  _RAND_373 = {1{`RANDOM}};
  cache_37_line_1 = _RAND_373[31:0];
  _RAND_374 = {1{`RANDOM}};
  cache_37_line_2 = _RAND_374[31:0];
  _RAND_375 = {1{`RANDOM}};
  cache_37_line_3 = _RAND_375[31:0];
  _RAND_376 = {1{`RANDOM}};
  cache_37_line_4 = _RAND_376[31:0];
  _RAND_377 = {1{`RANDOM}};
  cache_37_line_5 = _RAND_377[31:0];
  _RAND_378 = {1{`RANDOM}};
  cache_37_line_6 = _RAND_378[31:0];
  _RAND_379 = {1{`RANDOM}};
  cache_37_line_7 = _RAND_379[31:0];
  _RAND_380 = {1{`RANDOM}};
  cache_38_validBit = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  cache_38_tag = _RAND_381[4:0];
  _RAND_382 = {1{`RANDOM}};
  cache_38_line_0 = _RAND_382[31:0];
  _RAND_383 = {1{`RANDOM}};
  cache_38_line_1 = _RAND_383[31:0];
  _RAND_384 = {1{`RANDOM}};
  cache_38_line_2 = _RAND_384[31:0];
  _RAND_385 = {1{`RANDOM}};
  cache_38_line_3 = _RAND_385[31:0];
  _RAND_386 = {1{`RANDOM}};
  cache_38_line_4 = _RAND_386[31:0];
  _RAND_387 = {1{`RANDOM}};
  cache_38_line_5 = _RAND_387[31:0];
  _RAND_388 = {1{`RANDOM}};
  cache_38_line_6 = _RAND_388[31:0];
  _RAND_389 = {1{`RANDOM}};
  cache_38_line_7 = _RAND_389[31:0];
  _RAND_390 = {1{`RANDOM}};
  cache_39_validBit = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  cache_39_tag = _RAND_391[4:0];
  _RAND_392 = {1{`RANDOM}};
  cache_39_line_0 = _RAND_392[31:0];
  _RAND_393 = {1{`RANDOM}};
  cache_39_line_1 = _RAND_393[31:0];
  _RAND_394 = {1{`RANDOM}};
  cache_39_line_2 = _RAND_394[31:0];
  _RAND_395 = {1{`RANDOM}};
  cache_39_line_3 = _RAND_395[31:0];
  _RAND_396 = {1{`RANDOM}};
  cache_39_line_4 = _RAND_396[31:0];
  _RAND_397 = {1{`RANDOM}};
  cache_39_line_5 = _RAND_397[31:0];
  _RAND_398 = {1{`RANDOM}};
  cache_39_line_6 = _RAND_398[31:0];
  _RAND_399 = {1{`RANDOM}};
  cache_39_line_7 = _RAND_399[31:0];
  _RAND_400 = {1{`RANDOM}};
  cache_40_validBit = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  cache_40_tag = _RAND_401[4:0];
  _RAND_402 = {1{`RANDOM}};
  cache_40_line_0 = _RAND_402[31:0];
  _RAND_403 = {1{`RANDOM}};
  cache_40_line_1 = _RAND_403[31:0];
  _RAND_404 = {1{`RANDOM}};
  cache_40_line_2 = _RAND_404[31:0];
  _RAND_405 = {1{`RANDOM}};
  cache_40_line_3 = _RAND_405[31:0];
  _RAND_406 = {1{`RANDOM}};
  cache_40_line_4 = _RAND_406[31:0];
  _RAND_407 = {1{`RANDOM}};
  cache_40_line_5 = _RAND_407[31:0];
  _RAND_408 = {1{`RANDOM}};
  cache_40_line_6 = _RAND_408[31:0];
  _RAND_409 = {1{`RANDOM}};
  cache_40_line_7 = _RAND_409[31:0];
  _RAND_410 = {1{`RANDOM}};
  cache_41_validBit = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  cache_41_tag = _RAND_411[4:0];
  _RAND_412 = {1{`RANDOM}};
  cache_41_line_0 = _RAND_412[31:0];
  _RAND_413 = {1{`RANDOM}};
  cache_41_line_1 = _RAND_413[31:0];
  _RAND_414 = {1{`RANDOM}};
  cache_41_line_2 = _RAND_414[31:0];
  _RAND_415 = {1{`RANDOM}};
  cache_41_line_3 = _RAND_415[31:0];
  _RAND_416 = {1{`RANDOM}};
  cache_41_line_4 = _RAND_416[31:0];
  _RAND_417 = {1{`RANDOM}};
  cache_41_line_5 = _RAND_417[31:0];
  _RAND_418 = {1{`RANDOM}};
  cache_41_line_6 = _RAND_418[31:0];
  _RAND_419 = {1{`RANDOM}};
  cache_41_line_7 = _RAND_419[31:0];
  _RAND_420 = {1{`RANDOM}};
  cache_42_validBit = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  cache_42_tag = _RAND_421[4:0];
  _RAND_422 = {1{`RANDOM}};
  cache_42_line_0 = _RAND_422[31:0];
  _RAND_423 = {1{`RANDOM}};
  cache_42_line_1 = _RAND_423[31:0];
  _RAND_424 = {1{`RANDOM}};
  cache_42_line_2 = _RAND_424[31:0];
  _RAND_425 = {1{`RANDOM}};
  cache_42_line_3 = _RAND_425[31:0];
  _RAND_426 = {1{`RANDOM}};
  cache_42_line_4 = _RAND_426[31:0];
  _RAND_427 = {1{`RANDOM}};
  cache_42_line_5 = _RAND_427[31:0];
  _RAND_428 = {1{`RANDOM}};
  cache_42_line_6 = _RAND_428[31:0];
  _RAND_429 = {1{`RANDOM}};
  cache_42_line_7 = _RAND_429[31:0];
  _RAND_430 = {1{`RANDOM}};
  cache_43_validBit = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  cache_43_tag = _RAND_431[4:0];
  _RAND_432 = {1{`RANDOM}};
  cache_43_line_0 = _RAND_432[31:0];
  _RAND_433 = {1{`RANDOM}};
  cache_43_line_1 = _RAND_433[31:0];
  _RAND_434 = {1{`RANDOM}};
  cache_43_line_2 = _RAND_434[31:0];
  _RAND_435 = {1{`RANDOM}};
  cache_43_line_3 = _RAND_435[31:0];
  _RAND_436 = {1{`RANDOM}};
  cache_43_line_4 = _RAND_436[31:0];
  _RAND_437 = {1{`RANDOM}};
  cache_43_line_5 = _RAND_437[31:0];
  _RAND_438 = {1{`RANDOM}};
  cache_43_line_6 = _RAND_438[31:0];
  _RAND_439 = {1{`RANDOM}};
  cache_43_line_7 = _RAND_439[31:0];
  _RAND_440 = {1{`RANDOM}};
  cache_44_validBit = _RAND_440[0:0];
  _RAND_441 = {1{`RANDOM}};
  cache_44_tag = _RAND_441[4:0];
  _RAND_442 = {1{`RANDOM}};
  cache_44_line_0 = _RAND_442[31:0];
  _RAND_443 = {1{`RANDOM}};
  cache_44_line_1 = _RAND_443[31:0];
  _RAND_444 = {1{`RANDOM}};
  cache_44_line_2 = _RAND_444[31:0];
  _RAND_445 = {1{`RANDOM}};
  cache_44_line_3 = _RAND_445[31:0];
  _RAND_446 = {1{`RANDOM}};
  cache_44_line_4 = _RAND_446[31:0];
  _RAND_447 = {1{`RANDOM}};
  cache_44_line_5 = _RAND_447[31:0];
  _RAND_448 = {1{`RANDOM}};
  cache_44_line_6 = _RAND_448[31:0];
  _RAND_449 = {1{`RANDOM}};
  cache_44_line_7 = _RAND_449[31:0];
  _RAND_450 = {1{`RANDOM}};
  cache_45_validBit = _RAND_450[0:0];
  _RAND_451 = {1{`RANDOM}};
  cache_45_tag = _RAND_451[4:0];
  _RAND_452 = {1{`RANDOM}};
  cache_45_line_0 = _RAND_452[31:0];
  _RAND_453 = {1{`RANDOM}};
  cache_45_line_1 = _RAND_453[31:0];
  _RAND_454 = {1{`RANDOM}};
  cache_45_line_2 = _RAND_454[31:0];
  _RAND_455 = {1{`RANDOM}};
  cache_45_line_3 = _RAND_455[31:0];
  _RAND_456 = {1{`RANDOM}};
  cache_45_line_4 = _RAND_456[31:0];
  _RAND_457 = {1{`RANDOM}};
  cache_45_line_5 = _RAND_457[31:0];
  _RAND_458 = {1{`RANDOM}};
  cache_45_line_6 = _RAND_458[31:0];
  _RAND_459 = {1{`RANDOM}};
  cache_45_line_7 = _RAND_459[31:0];
  _RAND_460 = {1{`RANDOM}};
  cache_46_validBit = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  cache_46_tag = _RAND_461[4:0];
  _RAND_462 = {1{`RANDOM}};
  cache_46_line_0 = _RAND_462[31:0];
  _RAND_463 = {1{`RANDOM}};
  cache_46_line_1 = _RAND_463[31:0];
  _RAND_464 = {1{`RANDOM}};
  cache_46_line_2 = _RAND_464[31:0];
  _RAND_465 = {1{`RANDOM}};
  cache_46_line_3 = _RAND_465[31:0];
  _RAND_466 = {1{`RANDOM}};
  cache_46_line_4 = _RAND_466[31:0];
  _RAND_467 = {1{`RANDOM}};
  cache_46_line_5 = _RAND_467[31:0];
  _RAND_468 = {1{`RANDOM}};
  cache_46_line_6 = _RAND_468[31:0];
  _RAND_469 = {1{`RANDOM}};
  cache_46_line_7 = _RAND_469[31:0];
  _RAND_470 = {1{`RANDOM}};
  cache_47_validBit = _RAND_470[0:0];
  _RAND_471 = {1{`RANDOM}};
  cache_47_tag = _RAND_471[4:0];
  _RAND_472 = {1{`RANDOM}};
  cache_47_line_0 = _RAND_472[31:0];
  _RAND_473 = {1{`RANDOM}};
  cache_47_line_1 = _RAND_473[31:0];
  _RAND_474 = {1{`RANDOM}};
  cache_47_line_2 = _RAND_474[31:0];
  _RAND_475 = {1{`RANDOM}};
  cache_47_line_3 = _RAND_475[31:0];
  _RAND_476 = {1{`RANDOM}};
  cache_47_line_4 = _RAND_476[31:0];
  _RAND_477 = {1{`RANDOM}};
  cache_47_line_5 = _RAND_477[31:0];
  _RAND_478 = {1{`RANDOM}};
  cache_47_line_6 = _RAND_478[31:0];
  _RAND_479 = {1{`RANDOM}};
  cache_47_line_7 = _RAND_479[31:0];
  _RAND_480 = {1{`RANDOM}};
  cache_48_validBit = _RAND_480[0:0];
  _RAND_481 = {1{`RANDOM}};
  cache_48_tag = _RAND_481[4:0];
  _RAND_482 = {1{`RANDOM}};
  cache_48_line_0 = _RAND_482[31:0];
  _RAND_483 = {1{`RANDOM}};
  cache_48_line_1 = _RAND_483[31:0];
  _RAND_484 = {1{`RANDOM}};
  cache_48_line_2 = _RAND_484[31:0];
  _RAND_485 = {1{`RANDOM}};
  cache_48_line_3 = _RAND_485[31:0];
  _RAND_486 = {1{`RANDOM}};
  cache_48_line_4 = _RAND_486[31:0];
  _RAND_487 = {1{`RANDOM}};
  cache_48_line_5 = _RAND_487[31:0];
  _RAND_488 = {1{`RANDOM}};
  cache_48_line_6 = _RAND_488[31:0];
  _RAND_489 = {1{`RANDOM}};
  cache_48_line_7 = _RAND_489[31:0];
  _RAND_490 = {1{`RANDOM}};
  cache_49_validBit = _RAND_490[0:0];
  _RAND_491 = {1{`RANDOM}};
  cache_49_tag = _RAND_491[4:0];
  _RAND_492 = {1{`RANDOM}};
  cache_49_line_0 = _RAND_492[31:0];
  _RAND_493 = {1{`RANDOM}};
  cache_49_line_1 = _RAND_493[31:0];
  _RAND_494 = {1{`RANDOM}};
  cache_49_line_2 = _RAND_494[31:0];
  _RAND_495 = {1{`RANDOM}};
  cache_49_line_3 = _RAND_495[31:0];
  _RAND_496 = {1{`RANDOM}};
  cache_49_line_4 = _RAND_496[31:0];
  _RAND_497 = {1{`RANDOM}};
  cache_49_line_5 = _RAND_497[31:0];
  _RAND_498 = {1{`RANDOM}};
  cache_49_line_6 = _RAND_498[31:0];
  _RAND_499 = {1{`RANDOM}};
  cache_49_line_7 = _RAND_499[31:0];
  _RAND_500 = {1{`RANDOM}};
  cache_50_validBit = _RAND_500[0:0];
  _RAND_501 = {1{`RANDOM}};
  cache_50_tag = _RAND_501[4:0];
  _RAND_502 = {1{`RANDOM}};
  cache_50_line_0 = _RAND_502[31:0];
  _RAND_503 = {1{`RANDOM}};
  cache_50_line_1 = _RAND_503[31:0];
  _RAND_504 = {1{`RANDOM}};
  cache_50_line_2 = _RAND_504[31:0];
  _RAND_505 = {1{`RANDOM}};
  cache_50_line_3 = _RAND_505[31:0];
  _RAND_506 = {1{`RANDOM}};
  cache_50_line_4 = _RAND_506[31:0];
  _RAND_507 = {1{`RANDOM}};
  cache_50_line_5 = _RAND_507[31:0];
  _RAND_508 = {1{`RANDOM}};
  cache_50_line_6 = _RAND_508[31:0];
  _RAND_509 = {1{`RANDOM}};
  cache_50_line_7 = _RAND_509[31:0];
  _RAND_510 = {1{`RANDOM}};
  cache_51_validBit = _RAND_510[0:0];
  _RAND_511 = {1{`RANDOM}};
  cache_51_tag = _RAND_511[4:0];
  _RAND_512 = {1{`RANDOM}};
  cache_51_line_0 = _RAND_512[31:0];
  _RAND_513 = {1{`RANDOM}};
  cache_51_line_1 = _RAND_513[31:0];
  _RAND_514 = {1{`RANDOM}};
  cache_51_line_2 = _RAND_514[31:0];
  _RAND_515 = {1{`RANDOM}};
  cache_51_line_3 = _RAND_515[31:0];
  _RAND_516 = {1{`RANDOM}};
  cache_51_line_4 = _RAND_516[31:0];
  _RAND_517 = {1{`RANDOM}};
  cache_51_line_5 = _RAND_517[31:0];
  _RAND_518 = {1{`RANDOM}};
  cache_51_line_6 = _RAND_518[31:0];
  _RAND_519 = {1{`RANDOM}};
  cache_51_line_7 = _RAND_519[31:0];
  _RAND_520 = {1{`RANDOM}};
  cache_52_validBit = _RAND_520[0:0];
  _RAND_521 = {1{`RANDOM}};
  cache_52_tag = _RAND_521[4:0];
  _RAND_522 = {1{`RANDOM}};
  cache_52_line_0 = _RAND_522[31:0];
  _RAND_523 = {1{`RANDOM}};
  cache_52_line_1 = _RAND_523[31:0];
  _RAND_524 = {1{`RANDOM}};
  cache_52_line_2 = _RAND_524[31:0];
  _RAND_525 = {1{`RANDOM}};
  cache_52_line_3 = _RAND_525[31:0];
  _RAND_526 = {1{`RANDOM}};
  cache_52_line_4 = _RAND_526[31:0];
  _RAND_527 = {1{`RANDOM}};
  cache_52_line_5 = _RAND_527[31:0];
  _RAND_528 = {1{`RANDOM}};
  cache_52_line_6 = _RAND_528[31:0];
  _RAND_529 = {1{`RANDOM}};
  cache_52_line_7 = _RAND_529[31:0];
  _RAND_530 = {1{`RANDOM}};
  cache_53_validBit = _RAND_530[0:0];
  _RAND_531 = {1{`RANDOM}};
  cache_53_tag = _RAND_531[4:0];
  _RAND_532 = {1{`RANDOM}};
  cache_53_line_0 = _RAND_532[31:0];
  _RAND_533 = {1{`RANDOM}};
  cache_53_line_1 = _RAND_533[31:0];
  _RAND_534 = {1{`RANDOM}};
  cache_53_line_2 = _RAND_534[31:0];
  _RAND_535 = {1{`RANDOM}};
  cache_53_line_3 = _RAND_535[31:0];
  _RAND_536 = {1{`RANDOM}};
  cache_53_line_4 = _RAND_536[31:0];
  _RAND_537 = {1{`RANDOM}};
  cache_53_line_5 = _RAND_537[31:0];
  _RAND_538 = {1{`RANDOM}};
  cache_53_line_6 = _RAND_538[31:0];
  _RAND_539 = {1{`RANDOM}};
  cache_53_line_7 = _RAND_539[31:0];
  _RAND_540 = {1{`RANDOM}};
  cache_54_validBit = _RAND_540[0:0];
  _RAND_541 = {1{`RANDOM}};
  cache_54_tag = _RAND_541[4:0];
  _RAND_542 = {1{`RANDOM}};
  cache_54_line_0 = _RAND_542[31:0];
  _RAND_543 = {1{`RANDOM}};
  cache_54_line_1 = _RAND_543[31:0];
  _RAND_544 = {1{`RANDOM}};
  cache_54_line_2 = _RAND_544[31:0];
  _RAND_545 = {1{`RANDOM}};
  cache_54_line_3 = _RAND_545[31:0];
  _RAND_546 = {1{`RANDOM}};
  cache_54_line_4 = _RAND_546[31:0];
  _RAND_547 = {1{`RANDOM}};
  cache_54_line_5 = _RAND_547[31:0];
  _RAND_548 = {1{`RANDOM}};
  cache_54_line_6 = _RAND_548[31:0];
  _RAND_549 = {1{`RANDOM}};
  cache_54_line_7 = _RAND_549[31:0];
  _RAND_550 = {1{`RANDOM}};
  cache_55_validBit = _RAND_550[0:0];
  _RAND_551 = {1{`RANDOM}};
  cache_55_tag = _RAND_551[4:0];
  _RAND_552 = {1{`RANDOM}};
  cache_55_line_0 = _RAND_552[31:0];
  _RAND_553 = {1{`RANDOM}};
  cache_55_line_1 = _RAND_553[31:0];
  _RAND_554 = {1{`RANDOM}};
  cache_55_line_2 = _RAND_554[31:0];
  _RAND_555 = {1{`RANDOM}};
  cache_55_line_3 = _RAND_555[31:0];
  _RAND_556 = {1{`RANDOM}};
  cache_55_line_4 = _RAND_556[31:0];
  _RAND_557 = {1{`RANDOM}};
  cache_55_line_5 = _RAND_557[31:0];
  _RAND_558 = {1{`RANDOM}};
  cache_55_line_6 = _RAND_558[31:0];
  _RAND_559 = {1{`RANDOM}};
  cache_55_line_7 = _RAND_559[31:0];
  _RAND_560 = {1{`RANDOM}};
  cache_56_validBit = _RAND_560[0:0];
  _RAND_561 = {1{`RANDOM}};
  cache_56_tag = _RAND_561[4:0];
  _RAND_562 = {1{`RANDOM}};
  cache_56_line_0 = _RAND_562[31:0];
  _RAND_563 = {1{`RANDOM}};
  cache_56_line_1 = _RAND_563[31:0];
  _RAND_564 = {1{`RANDOM}};
  cache_56_line_2 = _RAND_564[31:0];
  _RAND_565 = {1{`RANDOM}};
  cache_56_line_3 = _RAND_565[31:0];
  _RAND_566 = {1{`RANDOM}};
  cache_56_line_4 = _RAND_566[31:0];
  _RAND_567 = {1{`RANDOM}};
  cache_56_line_5 = _RAND_567[31:0];
  _RAND_568 = {1{`RANDOM}};
  cache_56_line_6 = _RAND_568[31:0];
  _RAND_569 = {1{`RANDOM}};
  cache_56_line_7 = _RAND_569[31:0];
  _RAND_570 = {1{`RANDOM}};
  cache_57_validBit = _RAND_570[0:0];
  _RAND_571 = {1{`RANDOM}};
  cache_57_tag = _RAND_571[4:0];
  _RAND_572 = {1{`RANDOM}};
  cache_57_line_0 = _RAND_572[31:0];
  _RAND_573 = {1{`RANDOM}};
  cache_57_line_1 = _RAND_573[31:0];
  _RAND_574 = {1{`RANDOM}};
  cache_57_line_2 = _RAND_574[31:0];
  _RAND_575 = {1{`RANDOM}};
  cache_57_line_3 = _RAND_575[31:0];
  _RAND_576 = {1{`RANDOM}};
  cache_57_line_4 = _RAND_576[31:0];
  _RAND_577 = {1{`RANDOM}};
  cache_57_line_5 = _RAND_577[31:0];
  _RAND_578 = {1{`RANDOM}};
  cache_57_line_6 = _RAND_578[31:0];
  _RAND_579 = {1{`RANDOM}};
  cache_57_line_7 = _RAND_579[31:0];
  _RAND_580 = {1{`RANDOM}};
  cache_58_validBit = _RAND_580[0:0];
  _RAND_581 = {1{`RANDOM}};
  cache_58_tag = _RAND_581[4:0];
  _RAND_582 = {1{`RANDOM}};
  cache_58_line_0 = _RAND_582[31:0];
  _RAND_583 = {1{`RANDOM}};
  cache_58_line_1 = _RAND_583[31:0];
  _RAND_584 = {1{`RANDOM}};
  cache_58_line_2 = _RAND_584[31:0];
  _RAND_585 = {1{`RANDOM}};
  cache_58_line_3 = _RAND_585[31:0];
  _RAND_586 = {1{`RANDOM}};
  cache_58_line_4 = _RAND_586[31:0];
  _RAND_587 = {1{`RANDOM}};
  cache_58_line_5 = _RAND_587[31:0];
  _RAND_588 = {1{`RANDOM}};
  cache_58_line_6 = _RAND_588[31:0];
  _RAND_589 = {1{`RANDOM}};
  cache_58_line_7 = _RAND_589[31:0];
  _RAND_590 = {1{`RANDOM}};
  cache_59_validBit = _RAND_590[0:0];
  _RAND_591 = {1{`RANDOM}};
  cache_59_tag = _RAND_591[4:0];
  _RAND_592 = {1{`RANDOM}};
  cache_59_line_0 = _RAND_592[31:0];
  _RAND_593 = {1{`RANDOM}};
  cache_59_line_1 = _RAND_593[31:0];
  _RAND_594 = {1{`RANDOM}};
  cache_59_line_2 = _RAND_594[31:0];
  _RAND_595 = {1{`RANDOM}};
  cache_59_line_3 = _RAND_595[31:0];
  _RAND_596 = {1{`RANDOM}};
  cache_59_line_4 = _RAND_596[31:0];
  _RAND_597 = {1{`RANDOM}};
  cache_59_line_5 = _RAND_597[31:0];
  _RAND_598 = {1{`RANDOM}};
  cache_59_line_6 = _RAND_598[31:0];
  _RAND_599 = {1{`RANDOM}};
  cache_59_line_7 = _RAND_599[31:0];
  _RAND_600 = {1{`RANDOM}};
  cache_60_validBit = _RAND_600[0:0];
  _RAND_601 = {1{`RANDOM}};
  cache_60_tag = _RAND_601[4:0];
  _RAND_602 = {1{`RANDOM}};
  cache_60_line_0 = _RAND_602[31:0];
  _RAND_603 = {1{`RANDOM}};
  cache_60_line_1 = _RAND_603[31:0];
  _RAND_604 = {1{`RANDOM}};
  cache_60_line_2 = _RAND_604[31:0];
  _RAND_605 = {1{`RANDOM}};
  cache_60_line_3 = _RAND_605[31:0];
  _RAND_606 = {1{`RANDOM}};
  cache_60_line_4 = _RAND_606[31:0];
  _RAND_607 = {1{`RANDOM}};
  cache_60_line_5 = _RAND_607[31:0];
  _RAND_608 = {1{`RANDOM}};
  cache_60_line_6 = _RAND_608[31:0];
  _RAND_609 = {1{`RANDOM}};
  cache_60_line_7 = _RAND_609[31:0];
  _RAND_610 = {1{`RANDOM}};
  cache_61_validBit = _RAND_610[0:0];
  _RAND_611 = {1{`RANDOM}};
  cache_61_tag = _RAND_611[4:0];
  _RAND_612 = {1{`RANDOM}};
  cache_61_line_0 = _RAND_612[31:0];
  _RAND_613 = {1{`RANDOM}};
  cache_61_line_1 = _RAND_613[31:0];
  _RAND_614 = {1{`RANDOM}};
  cache_61_line_2 = _RAND_614[31:0];
  _RAND_615 = {1{`RANDOM}};
  cache_61_line_3 = _RAND_615[31:0];
  _RAND_616 = {1{`RANDOM}};
  cache_61_line_4 = _RAND_616[31:0];
  _RAND_617 = {1{`RANDOM}};
  cache_61_line_5 = _RAND_617[31:0];
  _RAND_618 = {1{`RANDOM}};
  cache_61_line_6 = _RAND_618[31:0];
  _RAND_619 = {1{`RANDOM}};
  cache_61_line_7 = _RAND_619[31:0];
  _RAND_620 = {1{`RANDOM}};
  cache_62_validBit = _RAND_620[0:0];
  _RAND_621 = {1{`RANDOM}};
  cache_62_tag = _RAND_621[4:0];
  _RAND_622 = {1{`RANDOM}};
  cache_62_line_0 = _RAND_622[31:0];
  _RAND_623 = {1{`RANDOM}};
  cache_62_line_1 = _RAND_623[31:0];
  _RAND_624 = {1{`RANDOM}};
  cache_62_line_2 = _RAND_624[31:0];
  _RAND_625 = {1{`RANDOM}};
  cache_62_line_3 = _RAND_625[31:0];
  _RAND_626 = {1{`RANDOM}};
  cache_62_line_4 = _RAND_626[31:0];
  _RAND_627 = {1{`RANDOM}};
  cache_62_line_5 = _RAND_627[31:0];
  _RAND_628 = {1{`RANDOM}};
  cache_62_line_6 = _RAND_628[31:0];
  _RAND_629 = {1{`RANDOM}};
  cache_62_line_7 = _RAND_629[31:0];
  _RAND_630 = {1{`RANDOM}};
  cache_63_validBit = _RAND_630[0:0];
  _RAND_631 = {1{`RANDOM}};
  cache_63_tag = _RAND_631[4:0];
  _RAND_632 = {1{`RANDOM}};
  cache_63_line_0 = _RAND_632[31:0];
  _RAND_633 = {1{`RANDOM}};
  cache_63_line_1 = _RAND_633[31:0];
  _RAND_634 = {1{`RANDOM}};
  cache_63_line_2 = _RAND_634[31:0];
  _RAND_635 = {1{`RANDOM}};
  cache_63_line_3 = _RAND_635[31:0];
  _RAND_636 = {1{`RANDOM}};
  cache_63_line_4 = _RAND_636[31:0];
  _RAND_637 = {1{`RANDOM}};
  cache_63_line_5 = _RAND_637[31:0];
  _RAND_638 = {1{`RANDOM}};
  cache_63_line_6 = _RAND_638[31:0];
  _RAND_639 = {1{`RANDOM}};
  cache_63_line_7 = _RAND_639[31:0];
  _RAND_640 = {8{`RANDOM}};
  dataBuffer = _RAND_640[255:0];
  _RAND_641 = {1{`RANDOM}};
  addrsBuffer = _RAND_641[15:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CacheControl(
  input   clock,
  input   reset,
  input   io_inMemRead,
  input   io_inMemWrite,
  input   io_hit,
  output  io_valid,
  output  io_cacheEn,
  output  io_blockWriteEn,
  output  io_outMemRead,
  output  io_outMemWrite,
  output  io_sel
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg  state; // @[CacheControl.scala 22:22]
  wire  _T_1 = ~state; // @[CacheControl.scala 35:21]
  wire  _GEN_2 = state ? 1'h0 : state; // @[CacheControl.scala 35:21 48:17 22:22]
  wire  _GEN_4 = ~state ? 1'h0 : state; // @[CacheControl.scala 35:21 38:23]
  wire  _GEN_5 = ~state | _GEN_2; // @[CacheControl.scala 35:21 41:17]
  wire  _GEN_7 = io_hit & io_inMemWrite; // @[CacheControl.scala 31:18 33:15 24:28]
  wire  _GEN_8 = io_hit ? 1'h0 : _T_1; // @[CacheControl.scala 31:18 25:31]
  wire  _GEN_9 = io_hit ? 1'h0 : _GEN_4; // @[CacheControl.scala 31:18 26:32]
  wire  _GEN_10 = io_hit ? state : _GEN_5; // @[CacheControl.scala 31:18 22:22]
  wire  _GEN_15 = (io_inMemRead | io_inMemWrite) & _GEN_10; // @[CacheControl.scala 30:38 59:11]
  assign io_valid = (io_inMemRead | io_inMemWrite) & io_hit; // @[CacheControl.scala 30:38 53:11]
  assign io_cacheEn = (io_inMemRead | io_inMemWrite) & _GEN_7; // @[CacheControl.scala 30:38 54:13]
  assign io_blockWriteEn = (io_inMemRead | io_inMemWrite) & _GEN_9; // @[CacheControl.scala 30:38 56:17]
  assign io_outMemRead = (io_inMemRead | io_inMemWrite) & _GEN_8; // @[CacheControl.scala 30:38 55:16]
  assign io_outMemWrite = (io_inMemRead | io_inMemWrite) & _GEN_9; // @[CacheControl.scala 30:38 56:17]
  assign io_sel = (io_inMemRead | io_inMemWrite) & _GEN_9; // @[CacheControl.scala 30:38 56:17]
  always @(posedge clock) begin
    if (reset) begin // @[CacheControl.scala 22:22]
      state <= 1'h0; // @[CacheControl.scala 22:22]
    end else begin
      state <= _GEN_15;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AddresSelector(
  input         io_sel,
  input  [10:0] io_addrs,
  input  [10:0] io_bufferAddrs,
  output [10:0] io_out
);
  assign io_out = io_sel ? io_bufferAddrs : io_addrs; // @[Cache.scala 128:16]
endmodule
module Cache(
  input          clock,
  input          reset,
  input          io_inMemRead,
  input          io_inMemWrite,
  input  [15:0]  io_addrs,
  input  [31:0]  io_cpuWriteData,
  output [31:0]  io_cpuReadData,
  input  [1:0]   io_storeType,
  output         io_valid,
  output [255:0] io_readBlock,
  input  [255:0] io_writeBlock,
  output         io_outMemRead,
  output         io_outMemWrite,
  output [10:0]  io_bufferAddrs
);
  wire  cache_clock; // @[Cache.scala 92:21]
  wire  cache_reset; // @[Cache.scala 92:21]
  wire [15:0] cache_io_addrs; // @[Cache.scala 92:21]
  wire [31:0] cache_io_cpuWriteData; // @[Cache.scala 92:21]
  wire [31:0] cache_io_cpuReadData; // @[Cache.scala 92:21]
  wire [1:0] cache_io_storeType; // @[Cache.scala 92:21]
  wire  cache_io_cpuWriteEn; // @[Cache.scala 92:21]
  wire [10:0] cache_io_bufferAddrs; // @[Cache.scala 92:21]
  wire [255:0] cache_io_readBlock; // @[Cache.scala 92:21]
  wire [255:0] cache_io_writeBlock; // @[Cache.scala 92:21]
  wire  cache_io_blockWriteEn; // @[Cache.scala 92:21]
  wire  cache_io_hit; // @[Cache.scala 92:21]
  wire  cacheControl_clock; // @[Cache.scala 93:28]
  wire  cacheControl_reset; // @[Cache.scala 93:28]
  wire  cacheControl_io_inMemRead; // @[Cache.scala 93:28]
  wire  cacheControl_io_inMemWrite; // @[Cache.scala 93:28]
  wire  cacheControl_io_hit; // @[Cache.scala 93:28]
  wire  cacheControl_io_valid; // @[Cache.scala 93:28]
  wire  cacheControl_io_cacheEn; // @[Cache.scala 93:28]
  wire  cacheControl_io_blockWriteEn; // @[Cache.scala 93:28]
  wire  cacheControl_io_outMemRead; // @[Cache.scala 93:28]
  wire  cacheControl_io_outMemWrite; // @[Cache.scala 93:28]
  wire  cacheControl_io_sel; // @[Cache.scala 93:28]
  wire  selector_io_sel; // @[Cache.scala 94:24]
  wire [10:0] selector_io_addrs; // @[Cache.scala 94:24]
  wire [10:0] selector_io_bufferAddrs; // @[Cache.scala 94:24]
  wire [10:0] selector_io_out; // @[Cache.scala 94:24]
  L1 cache ( // @[Cache.scala 92:21]
    .clock(cache_clock),
    .reset(cache_reset),
    .io_addrs(cache_io_addrs),
    .io_cpuWriteData(cache_io_cpuWriteData),
    .io_cpuReadData(cache_io_cpuReadData),
    .io_storeType(cache_io_storeType),
    .io_cpuWriteEn(cache_io_cpuWriteEn),
    .io_bufferAddrs(cache_io_bufferAddrs),
    .io_readBlock(cache_io_readBlock),
    .io_writeBlock(cache_io_writeBlock),
    .io_blockWriteEn(cache_io_blockWriteEn),
    .io_hit(cache_io_hit)
  );
  CacheControl cacheControl ( // @[Cache.scala 93:28]
    .clock(cacheControl_clock),
    .reset(cacheControl_reset),
    .io_inMemRead(cacheControl_io_inMemRead),
    .io_inMemWrite(cacheControl_io_inMemWrite),
    .io_hit(cacheControl_io_hit),
    .io_valid(cacheControl_io_valid),
    .io_cacheEn(cacheControl_io_cacheEn),
    .io_blockWriteEn(cacheControl_io_blockWriteEn),
    .io_outMemRead(cacheControl_io_outMemRead),
    .io_outMemWrite(cacheControl_io_outMemWrite),
    .io_sel(cacheControl_io_sel)
  );
  AddresSelector selector ( // @[Cache.scala 94:24]
    .io_sel(selector_io_sel),
    .io_addrs(selector_io_addrs),
    .io_bufferAddrs(selector_io_bufferAddrs),
    .io_out(selector_io_out)
  );
  assign io_cpuReadData = cache_io_cpuReadData; // @[Cache.scala 111:18]
  assign io_valid = cacheControl_io_valid; // @[Cache.scala 112:12]
  assign io_readBlock = cache_io_readBlock; // @[Cache.scala 113:16]
  assign io_outMemRead = cacheControl_io_outMemRead; // @[Cache.scala 114:17]
  assign io_outMemWrite = cacheControl_io_outMemWrite; // @[Cache.scala 115:18]
  assign io_bufferAddrs = selector_io_out; // @[Cache.scala 116:18]
  assign cache_clock = clock;
  assign cache_reset = reset;
  assign cache_io_addrs = io_addrs; // @[Cache.scala 96:18]
  assign cache_io_cpuWriteData = io_cpuWriteData; // @[Cache.scala 97:25]
  assign cache_io_storeType = io_storeType; // @[Cache.scala 98:22]
  assign cache_io_cpuWriteEn = cacheControl_io_cacheEn; // @[Cache.scala 99:23]
  assign cache_io_writeBlock = io_writeBlock; // @[Cache.scala 100:23]
  assign cache_io_blockWriteEn = cacheControl_io_blockWriteEn; // @[Cache.scala 101:25]
  assign cacheControl_clock = clock;
  assign cacheControl_reset = reset;
  assign cacheControl_io_inMemRead = io_inMemRead; // @[Cache.scala 103:29]
  assign cacheControl_io_inMemWrite = io_inMemWrite; // @[Cache.scala 104:30]
  assign cacheControl_io_hit = cache_io_hit; // @[Cache.scala 105:23]
  assign selector_io_sel = cacheControl_io_sel; // @[Cache.scala 107:19]
  assign selector_io_addrs = io_addrs[15:5]; // @[Cache.scala 108:32]
  assign selector_io_bufferAddrs = cache_io_bufferAddrs; // @[Cache.scala 109:27]
endmodule
module Processor(
  input          clock,
  input          reset,
  input  [31:0]  io_instr,
  input  [255:0] io_memReadBlock,
  output [10:0]  io_memAdrrs,
  output [8:0]   io_instrAddrs,
  output [255:0] io_memWriteBlock,
  output         io_memRead,
  output         io_memWrite
);
  wire  core_clock; // @[Processor.scala 19:20]
  wire  core_reset; // @[Processor.scala 19:20]
  wire [31:0] core_io_instr; // @[Processor.scala 19:20]
  wire [31:0] core_io_memReadData; // @[Processor.scala 19:20]
  wire  core_io_valid; // @[Processor.scala 19:20]
  wire [8:0] core_io_instrAddrs; // @[Processor.scala 19:20]
  wire [31:0] core_io_ALUOut; // @[Processor.scala 19:20]
  wire [31:0] core_io_memWriteData; // @[Processor.scala 19:20]
  wire  core_io_memRead; // @[Processor.scala 19:20]
  wire  core_io_memWrite; // @[Processor.scala 19:20]
  wire [1:0] core_io_storeType; // @[Processor.scala 19:20]
  wire  cacheCore_clock; // @[Processor.scala 20:25]
  wire  cacheCore_reset; // @[Processor.scala 20:25]
  wire  cacheCore_io_inMemRead; // @[Processor.scala 20:25]
  wire  cacheCore_io_inMemWrite; // @[Processor.scala 20:25]
  wire [15:0] cacheCore_io_addrs; // @[Processor.scala 20:25]
  wire [31:0] cacheCore_io_cpuWriteData; // @[Processor.scala 20:25]
  wire [31:0] cacheCore_io_cpuReadData; // @[Processor.scala 20:25]
  wire [1:0] cacheCore_io_storeType; // @[Processor.scala 20:25]
  wire  cacheCore_io_valid; // @[Processor.scala 20:25]
  wire [255:0] cacheCore_io_readBlock; // @[Processor.scala 20:25]
  wire [255:0] cacheCore_io_writeBlock; // @[Processor.scala 20:25]
  wire  cacheCore_io_outMemRead; // @[Processor.scala 20:25]
  wire  cacheCore_io_outMemWrite; // @[Processor.scala 20:25]
  wire [10:0] cacheCore_io_bufferAddrs; // @[Processor.scala 20:25]
  wire [31:0] _cacheCore_io_addrs_T = core_io_ALUOut; // @[Processor.scala 28:40]
  Core core ( // @[Processor.scala 19:20]
    .clock(core_clock),
    .reset(core_reset),
    .io_instr(core_io_instr),
    .io_memReadData(core_io_memReadData),
    .io_valid(core_io_valid),
    .io_instrAddrs(core_io_instrAddrs),
    .io_ALUOut(core_io_ALUOut),
    .io_memWriteData(core_io_memWriteData),
    .io_memRead(core_io_memRead),
    .io_memWrite(core_io_memWrite),
    .io_storeType(core_io_storeType)
  );
  Cache cacheCore ( // @[Processor.scala 20:25]
    .clock(cacheCore_clock),
    .reset(cacheCore_reset),
    .io_inMemRead(cacheCore_io_inMemRead),
    .io_inMemWrite(cacheCore_io_inMemWrite),
    .io_addrs(cacheCore_io_addrs),
    .io_cpuWriteData(cacheCore_io_cpuWriteData),
    .io_cpuReadData(cacheCore_io_cpuReadData),
    .io_storeType(cacheCore_io_storeType),
    .io_valid(cacheCore_io_valid),
    .io_readBlock(cacheCore_io_readBlock),
    .io_writeBlock(cacheCore_io_writeBlock),
    .io_outMemRead(cacheCore_io_outMemRead),
    .io_outMemWrite(cacheCore_io_outMemWrite),
    .io_bufferAddrs(cacheCore_io_bufferAddrs)
  );
  assign io_memAdrrs = cacheCore_io_bufferAddrs; // @[Processor.scala 37:15]
  assign io_instrAddrs = core_io_instrAddrs; // @[Processor.scala 33:17]
  assign io_memWriteBlock = cacheCore_io_readBlock; // @[Processor.scala 34:20]
  assign io_memRead = cacheCore_io_outMemRead; // @[Processor.scala 35:14]
  assign io_memWrite = cacheCore_io_outMemWrite; // @[Processor.scala 36:15]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_instr = io_instr; // @[Processor.scala 22:17]
  assign core_io_memReadData = cacheCore_io_cpuReadData; // @[Processor.scala 23:23]
  assign core_io_valid = cacheCore_io_valid; // @[Processor.scala 24:17]
  assign cacheCore_clock = clock;
  assign cacheCore_reset = reset;
  assign cacheCore_io_inMemRead = core_io_memRead; // @[Processor.scala 26:26]
  assign cacheCore_io_inMemWrite = core_io_memWrite; // @[Processor.scala 27:27]
  assign cacheCore_io_addrs = _cacheCore_io_addrs_T[15:0]; // @[Processor.scala 28:46]
  assign cacheCore_io_cpuWriteData = core_io_memWriteData; // @[Processor.scala 29:29]
  assign cacheCore_io_storeType = core_io_storeType; // @[Processor.scala 30:26]
  assign cacheCore_io_writeBlock = io_memReadBlock; // @[Processor.scala 31:27]
endmodule
